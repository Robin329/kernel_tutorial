// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.10.3.144
// Netlist written on Mon Nov 30 22:55:04 2020
//
// Verilog Description of module top
//

module top (clk_in, sw, key, seg_led_1, seg_led_2, rgb, led1, 
            led2, led3, led4, led5, led6, led7, led8) /* synthesis syn_module_defined=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(7[8:11])
    input clk_in;   // f:/home/mini-mcu/step_fpga/top.v(9[8:14])
    input [3:0]sw;   // f:/home/mini-mcu/step_fpga/top.v(11[14:16])
    input [3:0]key;   // f:/home/mini-mcu/step_fpga/top.v(12[14:17])
    output [8:0]seg_led_1;   // f:/home/mini-mcu/step_fpga/top.v(14[15:24])
    output [8:0]seg_led_2;   // f:/home/mini-mcu/step_fpga/top.v(15[15:24])
    output [2:0]rgb;   // f:/home/mini-mcu/step_fpga/top.v(17[17:20])
    output led1;   // f:/home/mini-mcu/step_fpga/top.v(19[9:13])
    output led2;   // f:/home/mini-mcu/step_fpga/top.v(20[9:13])
    output led3;   // f:/home/mini-mcu/step_fpga/top.v(21[9:13])
    output led4;   // f:/home/mini-mcu/step_fpga/top.v(22[9:13])
    output led5;   // f:/home/mini-mcu/step_fpga/top.v(23[9:13])
    output led6;   // f:/home/mini-mcu/step_fpga/top.v(24[9:13])
    output led7;   // f:/home/mini-mcu/step_fpga/top.v(25[9:13])
    output led8;   // f:/home/mini-mcu/step_fpga/top.v(26[9:13])
    
    wire clk_in_c /* synthesis SET_AS_NETWORK=clk_in_c, is_clock=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(9[8:14])
    wire [17:0]instruction /* synthesis syn_ramstyle="block_ram", ram_style="distributed" */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    
    wire GND_net, VCC_net, sw_c_3, sw_c_2, sw_c_1, sw_c_0, key_c_3, 
        key_c_2, key_c_1, key_c_0, seg_led_1_c_6, seg_led_1_c_5, seg_led_1_c_4, 
        seg_led_1_c_3, seg_led_1_c_2, seg_led_1_c_1, seg_led_1_c_0, 
        seg_led_2_c_6, seg_led_2_c_5, seg_led_2_c_4, seg_led_2_c_3, 
        seg_led_2_c_2, seg_led_2_c_1, seg_led_2_c_0, rgb_c_2, rgb_c_1, 
        rgb_c_0, led1_c_0, led2_c_1, led3_c_2, led4_c_3, led5_c_4, 
        led6_c_5, led7_c_6, led8_c_7, rst_n_in;
    wire [31:0]cnt;   // f:/home/mini-mcu/step_fpga/top.v(34[11:14])
    
    wire interrupt;
    wire [11:0]address;   // f:/home/mini-mcu/step_fpga/top.v(58[12:19])
    
    wire write_strobe;
    wire [7:0]in_port;   // f:/home/mini-mcu/step_fpga/top.v(61[11:18])
    wire [7:0]port_id;   // f:/home/mini-mcu/step_fpga/top.v(62[12:19])
    wire [7:0]out_port;   // f:/home/mini-mcu/step_fpga/top.v(62[21:29])
    wire [3:0]seg_data_1;   // f:/home/mini-mcu/step_fpga/top.v(64[10:20])
    wire [3:0]seg_data_2;   // f:/home/mini-mcu/step_fpga/top.v(64[22:32])
    
    wire cnt_31__N_88, rst_n_in_N_109, n14335, n153, n144, n857, 
        n156, n155, n154, n32, n150, n160, n14334, n10, in_port_7__N_37;
    wire [23:0]cnt_p;   // f:/home/mini-mcu/step_fpga/divide.v(27[22:27])
    
    wire n163, n14333, n158, n16312, n149, n143, n2071, n2075, 
        n2081, n2085, n142, n141, n8, n148, clk_in_c_enable_176, 
        n151, clk_in_c_enable_154, n147, n140, clk_in_c_enable_178, 
        n146, n139, n14332, n138, n16315, n16316, n16289, n16276, 
        n16290, n16277, n16351, n16348, n16260, n16261, n7942, 
        n7941, n7940, n7939, n16319, n80, n81, n82, n83, n16278, 
        n16279, n16330, n16264, n7934, n7933, n7932, n7931, n16336, 
        n114, n115, n116, n117, n7919, n7920, n7921, n7922, 
        n16346, n142_adj_1664, n143_adj_1665, n145, n146_adj_1666, 
        n16332, n16285, n16284, n16327, n16345, n16392, n7646, 
        n11714, n164, n165, n152, n162, n161, n137, n157, n31, 
        n1693, n136, n135, n134, n14331, n7, n8_adj_1667, n14330, 
        n14329, n159, n7_adj_1668, n10_adj_1669, n9, n145_adj_1670, 
        n14328, n9_adj_1671, n14327, n8_adj_1672, n14409, clk_in_c_enable_209, 
        n14326, n14302, n14325, n14324, n14301, n14323, n206, 
        n14322, n14300, n14299, n16318, n14298, n14297, n14296, 
        n14321, n14295, n14294, n14320, n14293, n14292, n14319, 
        n14318, n14317, n14316, n14315, n14291, n14290, n14289, 
        n14288, n14287, n11778, n7876, n7908, n16265, n7726, n7762, 
        n22301, n22297, n7623, n14339, n14338, n14337, n14336, 
        n16598, n14, n10_adj_1673, n16421, n16417, n22109;
    
    VHI i2 (.Z(VCC_net));
    \divide(N=12000000)  u1 (.interrupt(interrupt), .clk_in_c(clk_in_c), 
            .n22301(n22301), .n857(n857), .\cnt_p[22] (cnt_p[22]), .\cnt_p[23] (cnt_p[23]), 
            .GND_net(GND_net), .n14409(n14409)) /* synthesis syn_module_defined=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(51[3] 55[2])
    FD1S1I in_port_7__I_0_i1 (.D(sw_c_0), .CK(in_port_7__N_37), .CD(n22297), 
           .Q(in_port[0]));   // f:/home/mini-mcu/step_fpga/top.v(78[1] 85[4])
    defparam in_port_7__I_0_i1.GSR = "ENABLED";
    FD1P3AX out_i0_i6 (.D(out_port[5]), .SP(clk_in_c_enable_176), .CK(clk_in_c), 
            .Q(led6_c_5));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam out_i0_i6.GSR = "ENABLED";
    FD1P3AX rgb_i0_i1 (.D(out_port[0]), .SP(clk_in_c_enable_154), .CK(clk_in_c), 
            .Q(rgb_c_0));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam rgb_i0_i1.GSR = "ENABLED";
    FD1P3AX seg_data_2_i0_i0 (.D(out_port[0]), .SP(clk_in_c_enable_178), 
            .CK(clk_in_c), .Q(seg_data_2[0]));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam seg_data_2_i0_i0.GSR = "ENABLED";
    FD1S3JX rst_n_in_80 (.D(rst_n_in_N_109), .CK(clk_in_c), .PD(cnt_31__N_88), 
            .Q(rst_n_in));   // f:/home/mini-mcu/step_fpga/top.v(35[8] 46[4])
    defparam rst_n_in_80.GSR = "ENABLED";
    FD1S1I in_port_7__I_0_i2 (.D(sw_c_1), .CK(in_port_7__N_37), .CD(n22297), 
           .Q(in_port[1]));   // f:/home/mini-mcu/step_fpga/top.v(78[1] 85[4])
    defparam in_port_7__I_0_i2.GSR = "ENABLED";
    FD1S1I in_port_7__I_0_i3 (.D(sw_c_2), .CK(in_port_7__N_37), .CD(n22297), 
           .Q(in_port[2]));   // f:/home/mini-mcu/step_fpga/top.v(78[1] 85[4])
    defparam in_port_7__I_0_i3.GSR = "ENABLED";
    FD1S1I in_port_7__I_0_i4 (.D(sw_c_3), .CK(in_port_7__N_37), .CD(n22297), 
           .Q(in_port[3]));   // f:/home/mini-mcu/step_fpga/top.v(78[1] 85[4])
    defparam in_port_7__I_0_i4.GSR = "ENABLED";
    FD1S1I in_port_7__I_0_i5 (.D(key_c_0), .CK(in_port_7__N_37), .CD(n22297), 
           .Q(in_port[4]));   // f:/home/mini-mcu/step_fpga/top.v(78[1] 85[4])
    defparam in_port_7__I_0_i5.GSR = "ENABLED";
    FD1S1I in_port_7__I_0_i6 (.D(key_c_1), .CK(in_port_7__N_37), .CD(n22297), 
           .Q(in_port[5]));   // f:/home/mini-mcu/step_fpga/top.v(78[1] 85[4])
    defparam in_port_7__I_0_i6.GSR = "ENABLED";
    FD1S1I in_port_7__I_0_i7 (.D(key_c_2), .CK(in_port_7__N_37), .CD(n22297), 
           .Q(in_port[6]));   // f:/home/mini-mcu/step_fpga/top.v(78[1] 85[4])
    defparam in_port_7__I_0_i7.GSR = "ENABLED";
    FD1S1I in_port_7__I_0_i8 (.D(key_c_3), .CK(in_port_7__N_37), .CD(n22297), 
           .Q(in_port[7]));   // f:/home/mini-mcu/step_fpga/top.v(78[1] 85[4])
    defparam in_port_7__I_0_i8.GSR = "ENABLED";
    FD1P3AX out_i0_i5 (.D(out_port[4]), .SP(clk_in_c_enable_176), .CK(clk_in_c), 
            .Q(led5_c_4));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam out_i0_i5.GSR = "ENABLED";
    IB sw_pad_3 (.I(sw[3]), .O(sw_c_3));   // f:/home/mini-mcu/step_fpga/top.v(11[14:16])
    IB clk_in_pad (.I(clk_in), .O(clk_in_c));   // f:/home/mini-mcu/step_fpga/top.v(9[8:14])
    OB led8_pad (.I(led8_c_7), .O(led8));   // f:/home/mini-mcu/step_fpga/top.v(26[9:13])
    CCU2D cnt_830_add_4_15 (.A0(cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14293), .COUT(n14294), .S0(n152), .S1(n151));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_15.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_15.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_15.INJECT1_0 = "NO";
    defparam cnt_830_add_4_15.INJECT1_1 = "NO";
    CCU2D add_11182_2 (.A0(cnt[3]), .B0(cnt[2]), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n14326));
    defparam add_11182_2.INIT0 = 16'h1000;
    defparam add_11182_2.INIT1 = 16'h5555;
    defparam add_11182_2.INJECT1_0 = "NO";
    defparam add_11182_2.INJECT1_1 = "NO";
    CCU2D add_11181_24 (.A0(cnt[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14325), 
          .S1(cnt_31__N_88));
    defparam add_11181_24.INIT0 = 16'h5555;
    defparam add_11181_24.INIT1 = 16'h0000;
    defparam add_11181_24.INJECT1_0 = "NO";
    defparam add_11181_24.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_13 (.A0(cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14292), .COUT(n14293), .S0(n154), .S1(n153));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_13.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_13.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_13.INJECT1_0 = "NO";
    defparam cnt_830_add_4_13.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14291), 
          .COUT(n14292), .S0(n156), .S1(n155));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_11.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_11.INJECT1_0 = "NO";
    defparam cnt_830_add_4_11.INJECT1_1 = "NO";
    OB seg_led_1_pad_7 (.I(GND_net), .O(seg_led_1[7]));   // f:/home/mini-mcu/step_fpga/top.v(14[15:24])
    OB led7_pad (.I(led7_c_6), .O(led7));   // f:/home/mini-mcu/step_fpga/top.v(25[9:13])
    OB led6_pad (.I(led6_c_5), .O(led6));   // f:/home/mini-mcu/step_fpga/top.v(24[9:13])
    CCU2D cnt_830_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14290), 
          .COUT(n14291), .S0(n158), .S1(n157));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_9.INJECT1_0 = "NO";
    defparam cnt_830_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14289), 
          .COUT(n14290), .S0(n160), .S1(n159));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_7.INJECT1_0 = "NO";
    defparam cnt_830_add_4_7.INJECT1_1 = "NO";
    OB seg_led_1_pad_8 (.I(GND_net), .O(seg_led_1[8]));   // f:/home/mini-mcu/step_fpga/top.v(14[15:24])
    FD1P3AX out_i0_i4 (.D(out_port[3]), .SP(clk_in_c_enable_176), .CK(clk_in_c), 
            .Q(led4_c_3));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam out_i0_i4.GSR = "ENABLED";
    OB led5_pad (.I(led5_c_4), .O(led5));   // f:/home/mini-mcu/step_fpga/top.v(23[9:13])
    IB key_pad_0 (.I(key[0]), .O(key_c_0));   // f:/home/mini-mcu/step_fpga/top.v(12[14:17])
    CCU2D add_11181_22 (.A0(cnt[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14324), 
          .COUT(n14325));
    defparam add_11181_22.INIT0 = 16'h5555;
    defparam add_11181_22.INIT1 = 16'h5555;
    defparam add_11181_22.INJECT1_0 = "NO";
    defparam add_11181_22.INJECT1_1 = "NO";
    IB key_pad_1 (.I(key[1]), .O(key_c_1));   // f:/home/mini-mcu/step_fpga/top.v(12[14:17])
    FD1P3AX out_i0_i3 (.D(out_port[2]), .SP(clk_in_c_enable_176), .CK(clk_in_c), 
            .Q(led3_c_2));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam out_i0_i3.GSR = "ENABLED";
    IB key_pad_2 (.I(key[2]), .O(key_c_2));   // f:/home/mini-mcu/step_fpga/top.v(12[14:17])
    FD1P3AX seg_data_1_i0_i0 (.D(out_port[4]), .SP(clk_in_c_enable_178), 
            .CK(clk_in_c), .Q(seg_data_1[0]));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam seg_data_1_i0_i0.GSR = "ENABLED";
    IB key_pad_3 (.I(key[3]), .O(key_c_3));   // f:/home/mini-mcu/step_fpga/top.v(12[14:17])
    IB sw_pad_0 (.I(sw[0]), .O(sw_c_0));   // f:/home/mini-mcu/step_fpga/top.v(11[14:16])
    IB sw_pad_1 (.I(sw[1]), .O(sw_c_1));   // f:/home/mini-mcu/step_fpga/top.v(11[14:16])
    CCU2D add_11181_20 (.A0(cnt[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14323), 
          .COUT(n14324));
    defparam add_11181_20.INIT0 = 16'h5555;
    defparam add_11181_20.INIT1 = 16'h5555;
    defparam add_11181_20.INJECT1_0 = "NO";
    defparam add_11181_20.INJECT1_1 = "NO";
    IB sw_pad_2 (.I(sw[2]), .O(sw_c_2));   // f:/home/mini-mcu/step_fpga/top.v(11[14:16])
    CCU2D add_11181_18 (.A0(cnt[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14322), 
          .COUT(n14323));
    defparam add_11181_18.INIT0 = 16'h5555;
    defparam add_11181_18.INIT1 = 16'h5555;
    defparam add_11181_18.INJECT1_0 = "NO";
    defparam add_11181_18.INJECT1_1 = "NO";
    FD1P3AX out_i0_i2 (.D(out_port[1]), .SP(clk_in_c_enable_176), .CK(clk_in_c), 
            .Q(led2_c_1));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam out_i0_i2.GSR = "ENABLED";
    OB led4_pad (.I(led4_c_3), .O(led4));   // f:/home/mini-mcu/step_fpga/top.v(22[9:13])
    FD1P3AX out_i0_i1 (.D(out_port[0]), .SP(clk_in_c_enable_176), .CK(clk_in_c), 
            .Q(led1_c_0));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam out_i0_i1.GSR = "ENABLED";
    CCU2D cnt_830_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14288), 
          .COUT(n14289), .S0(n162), .S1(n161));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_5.INJECT1_0 = "NO";
    defparam cnt_830_add_4_5.INJECT1_1 = "NO";
    OB led3_pad (.I(led3_c_2), .O(led3));   // f:/home/mini-mcu/step_fpga/top.v(21[9:13])
    OB led2_pad (.I(led2_c_1), .O(led2));   // f:/home/mini-mcu/step_fpga/top.v(20[9:13])
    OB led1_pad (.I(led1_c_0), .O(led1));   // f:/home/mini-mcu/step_fpga/top.v(19[9:13])
    OB rgb_pad_0 (.I(rgb_c_0), .O(rgb[0]));   // f:/home/mini-mcu/step_fpga/top.v(17[17:20])
    OB rgb_pad_1 (.I(rgb_c_1), .O(rgb[1]));   // f:/home/mini-mcu/step_fpga/top.v(17[17:20])
    OB rgb_pad_2 (.I(rgb_c_2), .O(rgb[2]));   // f:/home/mini-mcu/step_fpga/top.v(17[17:20])
    OB seg_led_2_pad_0 (.I(seg_led_2_c_0), .O(seg_led_2[0]));   // f:/home/mini-mcu/step_fpga/top.v(15[15:24])
    OB seg_led_2_pad_1 (.I(seg_led_2_c_1), .O(seg_led_2[1]));   // f:/home/mini-mcu/step_fpga/top.v(15[15:24])
    OB seg_led_2_pad_2 (.I(seg_led_2_c_2), .O(seg_led_2[2]));   // f:/home/mini-mcu/step_fpga/top.v(15[15:24])
    OB seg_led_2_pad_3 (.I(seg_led_2_c_3), .O(seg_led_2[3]));   // f:/home/mini-mcu/step_fpga/top.v(15[15:24])
    OB seg_led_2_pad_4 (.I(seg_led_2_c_4), .O(seg_led_2[4]));   // f:/home/mini-mcu/step_fpga/top.v(15[15:24])
    OB seg_led_2_pad_5 (.I(seg_led_2_c_5), .O(seg_led_2[5]));   // f:/home/mini-mcu/step_fpga/top.v(15[15:24])
    OB seg_led_2_pad_6 (.I(seg_led_2_c_6), .O(seg_led_2[6]));   // f:/home/mini-mcu/step_fpga/top.v(15[15:24])
    OB seg_led_2_pad_7 (.I(GND_net), .O(seg_led_2[7]));   // f:/home/mini-mcu/step_fpga/top.v(15[15:24])
    OB seg_led_2_pad_8 (.I(GND_net), .O(seg_led_2[8]));   // f:/home/mini-mcu/step_fpga/top.v(15[15:24])
    OB seg_led_1_pad_0 (.I(seg_led_1_c_0), .O(seg_led_1[0]));   // f:/home/mini-mcu/step_fpga/top.v(14[15:24])
    OB seg_led_1_pad_1 (.I(seg_led_1_c_1), .O(seg_led_1[1]));   // f:/home/mini-mcu/step_fpga/top.v(14[15:24])
    OB seg_led_1_pad_2 (.I(seg_led_1_c_2), .O(seg_led_1[2]));   // f:/home/mini-mcu/step_fpga/top.v(14[15:24])
    OB seg_led_1_pad_3 (.I(seg_led_1_c_3), .O(seg_led_1[3]));   // f:/home/mini-mcu/step_fpga/top.v(14[15:24])
    OB seg_led_1_pad_4 (.I(seg_led_1_c_4), .O(seg_led_1[4]));   // f:/home/mini-mcu/step_fpga/top.v(14[15:24])
    OB seg_led_1_pad_5 (.I(seg_led_1_c_5), .O(seg_led_1[5]));   // f:/home/mini-mcu/step_fpga/top.v(14[15:24])
    CCU2D add_11181_16 (.A0(cnt[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14321), 
          .COUT(n14322));
    defparam add_11181_16.INIT0 = 16'h5aaa;
    defparam add_11181_16.INIT1 = 16'h5555;
    defparam add_11181_16.INJECT1_0 = "NO";
    defparam add_11181_16.INJECT1_1 = "NO";
    VLO i1 (.Z(GND_net));
    FD1P3AX cnt_830__i0 (.D(n165), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(n32)) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i0.GSR = "ENABLED";
    CCU2D add_11181_14 (.A0(cnt[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14320), 
          .COUT(n14321));
    defparam add_11181_14.INIT0 = 16'h5aaa;
    defparam add_11181_14.INIT1 = 16'h5555;
    defparam add_11181_14.INJECT1_0 = "NO";
    defparam add_11181_14.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_3 (.A0(n31), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14287), 
          .COUT(n14288), .S0(n164), .S1(n163));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_3.INJECT1_0 = "NO";
    defparam cnt_830_add_4_3.INJECT1_1 = "NO";
    FD1P3AX seg_data_2_i0_i3 (.D(out_port[3]), .SP(clk_in_c_enable_178), 
            .CK(clk_in_c), .Q(seg_data_2[3]));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam seg_data_2_i0_i3.GSR = "ENABLED";
    FD1P3AX seg_data_2_i0_i2 (.D(out_port[2]), .SP(clk_in_c_enable_178), 
            .CK(clk_in_c), .Q(seg_data_2[2]));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam seg_data_2_i0_i2.GSR = "ENABLED";
    FD1P3AX seg_data_2_i0_i1 (.D(out_port[1]), .SP(clk_in_c_enable_178), 
            .CK(clk_in_c), .Q(seg_data_2[1]));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam seg_data_2_i0_i1.GSR = "ENABLED";
    FD1P3AX rgb_i0_i3 (.D(out_port[2]), .SP(clk_in_c_enable_154), .CK(clk_in_c), 
            .Q(rgb_c_2));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam rgb_i0_i3.GSR = "ENABLED";
    FD1P3AX rgb_i0_i2 (.D(out_port[1]), .SP(clk_in_c_enable_154), .CK(clk_in_c), 
            .Q(rgb_c_1));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam rgb_i0_i2.GSR = "ENABLED";
    FD1P3AX out_i0_i8 (.D(out_port[7]), .SP(clk_in_c_enable_176), .CK(clk_in_c), 
            .Q(led8_c_7));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam out_i0_i8.GSR = "ENABLED";
    OB seg_led_1_pad_6 (.I(seg_led_1_c_6), .O(seg_led_1[6]));   // f:/home/mini-mcu/step_fpga/top.v(14[15:24])
    CCU2D cnt_830_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n32), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n14287), 
          .S1(n165));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_1.INIT0 = 16'hF000;
    defparam cnt_830_add_4_1.INIT1 = 16'h0555;
    defparam cnt_830_add_4_1.INJECT1_0 = "NO";
    defparam cnt_830_add_4_1.INJECT1_1 = "NO";
    CCU2D add_11181_12 (.A0(cnt[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14319), 
          .COUT(n14320));
    defparam add_11181_12.INIT0 = 16'h5555;
    defparam add_11181_12.INIT1 = 16'h5aaa;
    defparam add_11181_12.INJECT1_0 = "NO";
    defparam add_11181_12.INJECT1_1 = "NO";
    FD1P3AX seg_data_1_i0_i1 (.D(out_port[5]), .SP(clk_in_c_enable_178), 
            .CK(clk_in_c), .Q(seg_data_1[1]));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam seg_data_1_i0_i1.GSR = "ENABLED";
    CCU2D add_11181_10 (.A0(cnt[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14318), 
          .COUT(n14319));
    defparam add_11181_10.INIT0 = 16'h5aaa;
    defparam add_11181_10.INIT1 = 16'h5aaa;
    defparam add_11181_10.INJECT1_0 = "NO";
    defparam add_11181_10.INJECT1_1 = "NO";
    CCU2D add_11181_8 (.A0(cnt[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14317), 
          .COUT(n14318));
    defparam add_11181_8.INIT0 = 16'h5555;
    defparam add_11181_8.INIT1 = 16'h5aaa;
    defparam add_11181_8.INJECT1_0 = "NO";
    defparam add_11181_8.INJECT1_1 = "NO";
    FD1P3AX out_i0_i7 (.D(out_port[6]), .SP(clk_in_c_enable_176), .CK(clk_in_c), 
            .Q(led7_c_6));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam out_i0_i7.GSR = "ENABLED";
    GSR GSR_INST (.GSR(VCC_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 i2_3_lut (.A(port_id[0]), .B(port_id[1]), .C(n7623), .Z(clk_in_c_enable_154)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i2_3_lut.init = 16'h4040;
    LUT4 i6_4_lut (.A(port_id[3]), .B(port_id[1]), .C(port_id[5]), .D(port_id[7]), 
         .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/top.v(69[5:10])
    defparam i6_4_lut.init = 16'hfffe;
    FD1P3AX seg_data_1_i0_i2 (.D(out_port[6]), .SP(clk_in_c_enable_178), 
            .CK(clk_in_c), .Q(seg_data_1[2]));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam seg_data_1_i0_i2.GSR = "ENABLED";
    FD1P3AX seg_data_1_i0_i3 (.D(out_port[7]), .SP(clk_in_c_enable_178), 
            .CK(clk_in_c), .Q(seg_data_1[3]));   // f:/home/mini-mcu/step_fpga/top.v(66[8] 75[4])
    defparam seg_data_1_i0_i3.GSR = "ENABLED";
    FD1P3AX cnt_830__i1 (.D(n164), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(n31)) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i1.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(port_id[2]), .B(port_id[4]), .Z(n10_adj_1673)) /* synthesis lut_function=(A+(B)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(69[5:10])
    defparam i2_2_lut.init = 16'heeee;
    FD1P3AX cnt_830__i2 (.D(n163), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i2.GSR = "ENABLED";
    FD1P3AX cnt_830__i3 (.D(n162), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i3.GSR = "ENABLED";
    FD1P3AX cnt_830__i4 (.D(n161), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i4.GSR = "ENABLED";
    FD1P3AX cnt_830__i5 (.D(n160), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i5.GSR = "ENABLED";
    FD1P3AX cnt_830__i6 (.D(n159), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i6.GSR = "ENABLED";
    FD1P3AX cnt_830__i7 (.D(n158), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i7.GSR = "ENABLED";
    FD1P3AX cnt_830__i8 (.D(n157), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i8.GSR = "ENABLED";
    FD1P3AX cnt_830__i9 (.D(n156), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i9.GSR = "ENABLED";
    FD1P3AX cnt_830__i10 (.D(n155), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i10.GSR = "ENABLED";
    FD1P3AX cnt_830__i11 (.D(n154), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i11.GSR = "ENABLED";
    FD1P3AX cnt_830__i12 (.D(n153), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i12.GSR = "ENABLED";
    FD1P3AX cnt_830__i13 (.D(n152), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i13.GSR = "ENABLED";
    FD1P3AX cnt_830__i14 (.D(n151), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[14])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i14.GSR = "ENABLED";
    FD1P3AX cnt_830__i15 (.D(n150), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[15])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i15.GSR = "ENABLED";
    FD1P3AX cnt_830__i16 (.D(n149), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[16])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i16.GSR = "ENABLED";
    FD1P3AX cnt_830__i17 (.D(n148), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[17])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i17.GSR = "ENABLED";
    FD1P3AX cnt_830__i18 (.D(n147), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[18])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i18.GSR = "ENABLED";
    FD1P3AX cnt_830__i19 (.D(n146), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[19])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i19.GSR = "ENABLED";
    FD1P3AX cnt_830__i20 (.D(n145_adj_1670), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[20])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i20.GSR = "ENABLED";
    FD1P3AX cnt_830__i21 (.D(n144), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[21])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i21.GSR = "ENABLED";
    FD1P3AX cnt_830__i22 (.D(n143), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[22])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i22.GSR = "ENABLED";
    FD1P3AX cnt_830__i23 (.D(n142), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[23])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i23.GSR = "ENABLED";
    FD1P3AX cnt_830__i24 (.D(n141), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[24])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i24.GSR = "ENABLED";
    FD1P3AX cnt_830__i25 (.D(n140), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[25])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i25.GSR = "ENABLED";
    FD1P3AX cnt_830__i26 (.D(n139), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[26])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i26.GSR = "ENABLED";
    FD1P3AX cnt_830__i27 (.D(n138), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[27])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i27.GSR = "ENABLED";
    FD1P3AX cnt_830__i28 (.D(n137), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[28])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i28.GSR = "ENABLED";
    FD1P3AX cnt_830__i29 (.D(n136), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[29])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i29.GSR = "ENABLED";
    FD1P3AX cnt_830__i30 (.D(n135), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[30])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i30.GSR = "ENABLED";
    FD1P3AX cnt_830__i31 (.D(n134), .SP(clk_in_c_enable_209), .CK(clk_in_c), 
            .Q(cnt[31])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830__i31.GSR = "ENABLED";
    CCU2D add_11181_6 (.A0(cnt[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14316), 
          .COUT(n14317));
    defparam add_11181_6.INIT0 = 16'h5555;
    defparam add_11181_6.INIT1 = 16'h5555;
    defparam add_11181_6.INJECT1_0 = "NO";
    defparam add_11181_6.INJECT1_1 = "NO";
    CCU2D add_11181_4 (.A0(cnt[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14315), 
          .COUT(n14316));
    defparam add_11181_4.INIT0 = 16'h5aaa;
    defparam add_11181_4.INIT1 = 16'h5aaa;
    defparam add_11181_4.INJECT1_0 = "NO";
    defparam add_11181_4.INJECT1_1 = "NO";
    CCU2D add_11181_2 (.A0(cnt[9]), .B0(cnt[8]), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n14315));
    defparam add_11181_2.INIT0 = 16'h7000;
    defparam add_11181_2.INIT1 = 16'h5555;
    defparam add_11181_2.INJECT1_0 = "NO";
    defparam add_11181_2.INJECT1_1 = "NO";
    CCU2D add_11182_30 (.A0(cnt[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14339), 
          .S1(n1693));
    defparam add_11182_30.INIT0 = 16'h5555;
    defparam add_11182_30.INIT1 = 16'h0000;
    defparam add_11182_30.INJECT1_0 = "NO";
    defparam add_11182_30.INJECT1_1 = "NO";
    CCU2D add_11182_28 (.A0(cnt[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14338), 
          .COUT(n14339));
    defparam add_11182_28.INIT0 = 16'h5555;
    defparam add_11182_28.INIT1 = 16'h5555;
    defparam add_11182_28.INJECT1_0 = "NO";
    defparam add_11182_28.INJECT1_1 = "NO";
    CCU2D add_11182_26 (.A0(cnt[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14337), 
          .COUT(n14338));
    defparam add_11182_26.INIT0 = 16'h5555;
    defparam add_11182_26.INIT1 = 16'h5555;
    defparam add_11182_26.INJECT1_0 = "NO";
    defparam add_11182_26.INJECT1_1 = "NO";
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    CCU2D add_11182_24 (.A0(cnt[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14336), 
          .COUT(n14337));
    defparam add_11182_24.INIT0 = 16'h5555;
    defparam add_11182_24.INIT1 = 16'h5555;
    defparam add_11182_24.INJECT1_0 = "NO";
    defparam add_11182_24.INJECT1_1 = "NO";
    CCU2D add_11182_22 (.A0(cnt[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14335), 
          .COUT(n14336));
    defparam add_11182_22.INIT0 = 16'h5555;
    defparam add_11182_22.INIT1 = 16'h5555;
    defparam add_11182_22.INJECT1_0 = "NO";
    defparam add_11182_22.INJECT1_1 = "NO";
    LUT4 i6_4_lut_adj_268 (.A(port_id[3]), .B(n16598), .C(write_strobe), 
         .D(port_id[6]), .Z(n7623)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i6_4_lut_adj_268.init = 16'h0010;
    CCU2D add_11182_20 (.A0(cnt[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14334), 
          .COUT(n14335));
    defparam add_11182_20.INIT0 = 16'h5555;
    defparam add_11182_20.INIT1 = 16'h5555;
    defparam add_11182_20.INJECT1_0 = "NO";
    defparam add_11182_20.INJECT1_1 = "NO";
    rom rom (.address({address}), .clk_in_c(clk_in_c), .GND_net(GND_net), 
        .VCC_net(VCC_net), .instruction({instruction}), .n16312(n16312), 
        .n11778(n11778), .n16351(n16351), .n11714(n11714), .n16261(n16261), 
        .n7908(n7908), .n16392(n16392), .n7941(n7941), .n7762(n7762), 
        .n7726(n7726), .n82(n82), .n81(n81), .n7876(n7876), .n16315(n16315), 
        .n16417(n16417), .n22109(n22109), .n7646(n7646), .n2075(n2075), 
        .n9(n9), .n10(n10), .n8(n8), .n7(n7_adj_1668), .n83(n83), 
        .n7940(n7940), .n7942(n7942), .n2081(n2081), .n16348(n16348), 
        .n9_adj_6(n9_adj_1671), .n10_adj_7(n10_adj_1669), .n7_adj_8(n7), 
        .n8_adj_9(n8_adj_1667), .n16277(n16277), .n7939(n7939), .n16289(n16289), 
        .n7921(n7921), .n16345(n16345), .n7919(n7919), .n16285(n16285), 
        .n16332(n16332), .n145(n145), .n16284(n16284), .n16327(n16327), 
        .n7920(n7920), .n143(n143_adj_1665), .n142(n142_adj_1664), .n16290(n16290), 
        .n16346(n16346), .n7922(n7922), .n146(n146_adj_1666), .n2071(n2071), 
        .n8_adj_10(n8_adj_1672), .n16316(n16316), .n16260(n16260), .n2085(n2085), 
        .n206(n206), .n116(n116), .n16319(n16319), .n7934(n7934), .n16279(n16279), 
        .n7932(n7932), .n114(n114), .n16318(n16318), .n16278(n16278), 
        .n16330(n16330), .n115(n115), .n7933(n7933), .n16276(n16276), 
        .n80(n80), .n16264(n16264), .n16336(n16336), .n7931(n7931), 
        .n16265(n16265), .n117(n117), .n16421(n16421)) /* synthesis syn_module_defined=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(104[5] 109[2])
    LUT4 i6366_1_lut (.A(cnt_31__N_88), .Z(clk_in_c_enable_209)) /* synthesis lut_function=(!(A)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(34[11:14])
    defparam i6366_1_lut.init = 16'h5555;
    LUT4 i13430_4_lut (.A(port_id[7]), .B(port_id[5]), .C(port_id[2]), 
         .D(port_id[4]), .Z(n16598)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13430_4_lut.init = 16'hfffe;
    seg_display seg_display (.seg_data_1({seg_data_1}), .seg_led_1_c_5(seg_led_1_c_5), 
            .seg_led_1_c_6(seg_led_1_c_6), .seg_led_1_c_1(seg_led_1_c_1), 
            .seg_led_1_c_2(seg_led_1_c_2), .seg_led_1_c_3(seg_led_1_c_3), 
            .seg_data_2({seg_data_2}), .seg_led_2_c_2(seg_led_2_c_2), .seg_led_2_c_5(seg_led_2_c_5), 
            .seg_led_2_c_6(seg_led_2_c_6), .seg_led_2_c_1(seg_led_2_c_1), 
            .seg_led_2_c_3(seg_led_2_c_3), .seg_led_2_c_0(seg_led_2_c_0), 
            .seg_led_2_c_4(seg_led_2_c_4), .seg_led_1_c_0(seg_led_1_c_0), 
            .seg_led_1_c_4(seg_led_1_c_4)) /* synthesis syn_module_defined=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(113[13] 118[2])
    CCU2D add_11182_18 (.A0(cnt[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14333), 
          .COUT(n14334));
    defparam add_11182_18.INIT0 = 16'h5555;
    defparam add_11182_18.INIT1 = 16'h5555;
    defparam add_11182_18.INJECT1_0 = "NO";
    defparam add_11182_18.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut (.A(n7623), .B(port_id[1]), .C(port_id[0]), .Z(clk_in_c_enable_176)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_269 (.A(n7623), .B(port_id[1]), .C(port_id[0]), 
         .Z(clk_in_c_enable_178)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_269.init = 16'h0202;
    CCU2D add_11182_16 (.A0(cnt[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14332), 
          .COUT(n14333));
    defparam add_11182_16.INIT0 = 16'h5555;
    defparam add_11182_16.INIT1 = 16'h5555;
    defparam add_11182_16.INJECT1_0 = "NO";
    defparam add_11182_16.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_33 (.A0(cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14302), .S0(n134));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_33.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_33.INIT1 = 16'h0000;
    defparam cnt_830_add_4_33.INJECT1_0 = "NO";
    defparam cnt_830_add_4_33.INJECT1_1 = "NO";
    CCU2D add_11182_14 (.A0(cnt[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14331), 
          .COUT(n14332));
    defparam add_11182_14.INIT0 = 16'h5555;
    defparam add_11182_14.INIT1 = 16'h5555;
    defparam add_11182_14.INJECT1_0 = "NO";
    defparam add_11182_14.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_31 (.A0(cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14301), .COUT(n14302), .S0(n136), .S1(n135));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_31.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_31.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_31.INJECT1_0 = "NO";
    defparam cnt_830_add_4_31.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_29 (.A0(cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14300), .COUT(n14301), .S0(n138), .S1(n137));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_29.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_29.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_29.INJECT1_0 = "NO";
    defparam cnt_830_add_4_29.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_27 (.A0(cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14299), .COUT(n14300), .S0(n140), .S1(n139));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_27.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_27.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_27.INJECT1_0 = "NO";
    defparam cnt_830_add_4_27.INJECT1_1 = "NO";
    CCU2D add_11182_12 (.A0(cnt[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14330), 
          .COUT(n14331));
    defparam add_11182_12.INIT0 = 16'h5555;
    defparam add_11182_12.INIT1 = 16'h5555;
    defparam add_11182_12.INJECT1_0 = "NO";
    defparam add_11182_12.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_25 (.A0(cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14298), .COUT(n14299), .S0(n142), .S1(n141));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_25.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_25.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_25.INJECT1_0 = "NO";
    defparam cnt_830_add_4_25.INJECT1_1 = "NO";
    CCU2D add_11182_10 (.A0(cnt[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14329), 
          .COUT(n14330));
    defparam add_11182_10.INIT0 = 16'h5555;
    defparam add_11182_10.INIT1 = 16'h5555;
    defparam add_11182_10.INJECT1_0 = "NO";
    defparam add_11182_10.INJECT1_1 = "NO";
    CCU2D add_11182_8 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14328), 
          .COUT(n14329));
    defparam add_11182_8.INIT0 = 16'h5555;
    defparam add_11182_8.INIT1 = 16'h5555;
    defparam add_11182_8.INJECT1_0 = "NO";
    defparam add_11182_8.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_23 (.A0(cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14297), .COUT(n14298), .S0(n144), .S1(n143));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_23.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_23.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_23.INJECT1_0 = "NO";
    defparam cnt_830_add_4_23.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_21 (.A0(cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14296), .COUT(n14297), .S0(n146), .S1(n145_adj_1670));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_21.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_21.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_21.INJECT1_0 = "NO";
    defparam cnt_830_add_4_21.INJECT1_1 = "NO";
    CCU2D add_11182_6 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14327), 
          .COUT(n14328));
    defparam add_11182_6.INIT0 = 16'h5555;
    defparam add_11182_6.INIT1 = 16'h5555;
    defparam add_11182_6.INJECT1_0 = "NO";
    defparam add_11182_6.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_19 (.A0(cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14295), .COUT(n14296), .S0(n148), .S1(n147));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_19.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_19.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_19.INJECT1_0 = "NO";
    defparam cnt_830_add_4_19.INJECT1_1 = "NO";
    CCU2D add_11182_4 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14326), 
          .COUT(n14327));
    defparam add_11182_4.INIT0 = 16'h5aaa;
    defparam add_11182_4.INIT1 = 16'h5aaa;
    defparam add_11182_4.INJECT1_0 = "NO";
    defparam add_11182_4.INJECT1_1 = "NO";
    CCU2D cnt_830_add_4_17 (.A0(cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14294), .COUT(n14295), .S0(n150), .S1(n149));   // f:/home/mini-mcu/step_fpga/top.v(43[14:20])
    defparam cnt_830_add_4_17.INIT0 = 16'hfaaa;
    defparam cnt_830_add_4_17.INIT1 = 16'hfaaa;
    defparam cnt_830_add_4_17.INJECT1_0 = "NO";
    defparam cnt_830_add_4_17.INJECT1_1 = "NO";
    LUT4 i599_1_lut (.A(n1693), .Z(rst_n_in_N_109)) /* synthesis lut_function=(!(A)) */ ;
    defparam i599_1_lut.init = 16'h5555;
    LUT4 i7_4_lut_rep_730 (.A(port_id[0]), .B(n14), .C(n10_adj_1673), 
         .D(port_id[6]), .Z(n22297)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/top.v(69[5:10])
    defparam i7_4_lut_rep_730.init = 16'hfffe;
    LUT4 port_id_7__I_0_i16_1_lut_4_lut (.A(port_id[0]), .B(n14), .C(n10_adj_1673), 
         .D(port_id[6]), .Z(in_port_7__N_37)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/top.v(69[5:10])
    defparam port_id_7__I_0_i16_1_lut_4_lut.init = 16'h0001;
    mcu mcu (.clk_in_c(clk_in_c), .n11714(n11714), .instruction({instruction}), 
        .n22301(n22301), .interrupt(interrupt), .n16290(n16290), .out_port({out_port}), 
        .port_id({port_id}), .write_strobe(write_strobe), .GND_net(GND_net), 
        .address({address}), .VCC_net(VCC_net), .n7762(n7762), .n7908(n7908), 
        .n11778(n11778), .n16278(n16278), .n7876(n7876), .n16417(n16417), 
        .n16279(n16279), .n206(n206), .n7646(n7646), .n16312(n16312), 
        .n16392(n16392), .n22109(n22109), .n2085(n2085), .n7921(n7921), 
        .n2071(n2071), .n2081(n2081), .n7920(n7920), .n7726(n7726), 
        .n7919(n7919), .n16261(n16261), .n16284(n16284), .n2075(n2075), 
        .n16277(n16277), .n16260(n16260), .n16285(n16285), .n16276(n16276), 
        .n83(n83), .n146(n146_adj_1666), .n16421(n16421), .n82(n82), 
        .n81(n81), .n143(n143_adj_1665), .n80(n80), .n16351(n16351), 
        .n16327(n16327), .n16316(n16316), .n16348(n16348), .n16332(n16332), 
        .rst_n_in(rst_n_in), .n16315(n16315), .n7939(n7939), .n7922(n7922), 
        .n7940(n7940), .n7941(n7941), .n7942(n7942), .n9(n9_adj_1671), 
        .n9_adj_1(n9), .in_port({in_port}), .n7(n7), .n7_adj_2(n7_adj_1668), 
        .n10(n10_adj_1669), .n10_adj_3(n10), .n7931(n7931), .n8(n8_adj_1667), 
        .n8_adj_4(n8), .n16330(n16330), .n16336(n16336), .n115(n115), 
        .n117(n117), .n16264(n16264), .n16265(n16265), .n7934(n7934), 
        .n8_adj_5(n8_adj_1672), .n7933(n7933), .n7932(n7932), .\cnt_p[22] (cnt_p[22]), 
        .\cnt_p[23] (cnt_p[23]), .n14409(n14409), .n857(n857), .n16289(n16289), 
        .n16318(n16318), .n16319(n16319), .n114(n114), .n116(n116), 
        .n145(n145), .n142(n142_adj_1664), .n16346(n16346), .n16345(n16345)) /* synthesis syn_module_defined=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(90[5] 102[2])
    
endmodule
//
// Verilog Description of module \divide(N=12000000) 
//

module \divide(N=12000000)  (interrupt, clk_in_c, n22301, n857, \cnt_p[22] , 
            \cnt_p[23] , GND_net, n14409) /* synthesis syn_module_defined=1 */ ;
    output interrupt;
    input clk_in_c;
    input n22301;
    input n857;
    output \cnt_p[22] ;
    output \cnt_p[23] ;
    input GND_net;
    output n14409;
    
    wire clk_in_c /* synthesis SET_AS_NETWORK=clk_in_c, is_clock=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(9[8:14])
    
    wire clkout_N_161;
    wire [23:0]cnt_p;   // f:/home/mini-mcu/step_fpga/divide.v(27[22:27])
    wire [23:0]n101;
    
    wire n14314, n14313, n14312, n14311, n14310, n14309, n14308, 
        n14307, n14306, n14305, n14304, n14303, n14373, n16388, 
        n16386, n16478, n4, n12064, n16387, n4_adj_1663, n22, 
        n14348, n14, n10;
    
    FD1S3IX clk_p_29 (.D(clkout_N_161), .CK(clk_in_c), .CD(n22301), .Q(interrupt));   // f:/home/mini-mcu/step_fpga/divide.v(42[12] 50[6])
    defparam clk_p_29.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i0 (.D(n101[0]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[0])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i0.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i1 (.D(n101[1]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[1])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i1.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i2 (.D(n101[2]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[2])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i2.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i3 (.D(n101[3]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[3])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i3.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i4 (.D(n101[4]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[4])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i4.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i5 (.D(n101[5]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[5])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i5.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i6 (.D(n101[6]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[6])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i6.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i7 (.D(n101[7]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[7])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i7.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i8 (.D(n101[8]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[8])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i8.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i9 (.D(n101[9]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[9])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i9.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i10 (.D(n101[10]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[10])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i10.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i11 (.D(n101[11]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[11])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i11.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i12 (.D(n101[12]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[12])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i12.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i13 (.D(n101[13]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[13])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i13.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i14 (.D(n101[14]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[14])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i14.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i15 (.D(n101[15]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[15])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i15.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i16 (.D(n101[16]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[16])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i16.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i17 (.D(n101[17]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[17])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i17.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i18 (.D(n101[18]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[18])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i18.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i19 (.D(n101[19]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[19])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i19.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i20 (.D(n101[20]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[20])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i20.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i21 (.D(n101[21]), .CK(clk_in_c), .CD(n857), .Q(cnt_p[21])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i21.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i22 (.D(n101[22]), .CK(clk_in_c), .CD(n857), .Q(\cnt_p[22] )) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i22.GSR = "ENABLED";
    FD1S3IX cnt_p_831__i23 (.D(n101[23]), .CK(clk_in_c), .CD(n857), .Q(\cnt_p[23] )) /* synthesis syn_use_carry_chain=1 */ ;   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831__i23.GSR = "ENABLED";
    CCU2D cnt_p_831_add_4_25 (.A0(\cnt_p[23] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14314), .S0(n101[23]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_25.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_25.INIT1 = 16'h0000;
    defparam cnt_p_831_add_4_25.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_25.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_23 (.A0(cnt_p[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\cnt_p[22] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14313), .COUT(n14314), .S0(n101[21]), 
          .S1(n101[22]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_23.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_23.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_23.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_23.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_21 (.A0(cnt_p[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14312), .COUT(n14313), .S0(n101[19]), 
          .S1(n101[20]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_21.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_21.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_21.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_21.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_19 (.A0(cnt_p[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14311), .COUT(n14312), .S0(n101[17]), 
          .S1(n101[18]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_19.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_19.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_19.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_19.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_17 (.A0(cnt_p[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14310), .COUT(n14311), .S0(n101[15]), 
          .S1(n101[16]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_17.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_17.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_17.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_17.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_15 (.A0(cnt_p[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14309), .COUT(n14310), .S0(n101[13]), 
          .S1(n101[14]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_15.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_15.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_15.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_15.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_13 (.A0(cnt_p[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14308), .COUT(n14309), .S0(n101[11]), 
          .S1(n101[12]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_13.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_13.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_13.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_13.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_11 (.A0(cnt_p[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14307), .COUT(n14308), .S0(n101[9]), .S1(n101[10]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_11.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_11.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_9 (.A0(cnt_p[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14306), .COUT(n14307), .S0(n101[7]), .S1(n101[8]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_9.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_7 (.A0(cnt_p[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14305), .COUT(n14306), .S0(n101[5]), .S1(n101[6]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_7.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_5 (.A0(cnt_p[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14304), .COUT(n14305), .S0(n101[3]), .S1(n101[4]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_5.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_3 (.A0(cnt_p[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14303), .COUT(n14304), .S0(n101[1]), .S1(n101[2]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_p_831_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_p_831_add_4_3.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_p_831_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_p[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n14303), .S1(n101[0]));   // f:/home/mini-mcu/step_fpga/divide.v(38[16:23])
    defparam cnt_p_831_add_4_1.INIT0 = 16'hF000;
    defparam cnt_p_831_add_4_1.INIT1 = 16'h0555;
    defparam cnt_p_831_add_4_1.INJECT1_0 = "NO";
    defparam cnt_p_831_add_4_1.INJECT1_1 = "NO";
    LUT4 i9063_4_lut (.A(n14373), .B(\cnt_p[23] ), .C(\cnt_p[22] ), .D(cnt_p[21]), 
         .Z(clkout_N_161)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i9063_4_lut.init = 16'hfcec;
    LUT4 i2_4_lut (.A(cnt_p[20]), .B(n16388), .C(cnt_p[19]), .D(cnt_p[18]), 
         .Z(n14373)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'ha080;
    LUT4 i2_4_lut_adj_263 (.A(n16386), .B(n16478), .C(cnt_p[15]), .D(n4), 
         .Z(n16388)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_263.init = 16'ha080;
    LUT4 i1_4_lut (.A(cnt_p[11]), .B(cnt_p[12]), .C(n12064), .D(cnt_p[10]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'heccc;
    LUT4 i8925_3_lut (.A(cnt_p[7]), .B(cnt_p[9]), .C(cnt_p[8]), .Z(n12064)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i8925_3_lut.init = 16'hecec;
    LUT4 i1_2_lut (.A(cnt_p[17]), .B(cnt_p[16]), .Z(n16386)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_264 (.A(cnt_p[14]), .B(cnt_p[13]), .Z(n16478)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_264.init = 16'heeee;
    LUT4 i2_4_lut_adj_265 (.A(cnt_p[21]), .B(cnt_p[20]), .C(n16387), .D(cnt_p[19]), 
         .Z(n14409)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_265.init = 16'h8880;
    LUT4 i2_4_lut_adj_266 (.A(n16386), .B(n16478), .C(cnt_p[18]), .D(n4_adj_1663), 
         .Z(n16387)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_266.init = 16'ha080;
    LUT4 i1_4_lut_adj_267 (.A(cnt_p[12]), .B(cnt_p[15]), .C(cnt_p[11]), 
         .D(n22), .Z(n4_adj_1663)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_267.init = 16'heccc;
    LUT4 i970_4_lut (.A(n14348), .B(cnt_p[10]), .C(cnt_p[9]), .D(cnt_p[8]), 
         .Z(n22)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i970_4_lut.init = 16'hfcec;
    LUT4 i7_4_lut (.A(cnt_p[0]), .B(n14), .C(n10), .D(cnt_p[4]), .Z(n14348)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cnt_p[2]), .B(cnt_p[5]), .C(cnt_p[3]), .D(cnt_p[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i2_2_lut (.A(cnt_p[6]), .B(cnt_p[7]), .Z(n10)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module rom
//

module rom (address, clk_in_c, GND_net, VCC_net, instruction, n16312, 
            n11778, n16351, n11714, n16261, n7908, n16392, n7941, 
            n7762, n7726, n82, n81, n7876, n16315, n16417, n22109, 
            n7646, n2075, n9, n10, n8, n7, n83, n7940, n7942, 
            n2081, n16348, n9_adj_6, n10_adj_7, n7_adj_8, n8_adj_9, 
            n16277, n7939, n16289, n7921, n16345, n7919, n16285, 
            n16332, n145, n16284, n16327, n7920, n143, n142, n16290, 
            n16346, n7922, n146, n2071, n8_adj_10, n16316, n16260, 
            n2085, n206, n116, n16319, n7934, n16279, n7932, n114, 
            n16318, n16278, n16330, n115, n7933, n16276, n80, 
            n16264, n16336, n7931, n16265, n117, n16421) /* synthesis syn_module_defined=1 */ ;
    input [11:0]address;
    input clk_in_c;
    input GND_net;
    input VCC_net;
    output [17:0]instruction;
    input n16312;
    input n11778;
    output n16351;
    input n11714;
    output n16261;
    input n7908;
    input n16392;
    output n7941;
    input n7762;
    input n7726;
    output n82;
    output n81;
    input n7876;
    output n16315;
    output n16417;
    output n22109;
    input n7646;
    output n2075;
    output n9;
    output n10;
    output n8;
    output n7;
    output n83;
    output n7940;
    output n7942;
    output n2081;
    output n16348;
    output n9_adj_6;
    output n10_adj_7;
    output n7_adj_8;
    output n8_adj_9;
    output n16277;
    output n7939;
    output n16289;
    output n7921;
    output n16345;
    output n7919;
    output n16285;
    output n16332;
    output n145;
    output n16284;
    output n16327;
    output n7920;
    output n143;
    output n142;
    output n16290;
    output n16346;
    output n7922;
    output n146;
    output n2071;
    output n8_adj_10;
    output n16316;
    output n16260;
    output n2085;
    input n206;
    output n116;
    output n16319;
    output n7934;
    output n16279;
    output n7932;
    output n114;
    output n16318;
    output n16278;
    output n16330;
    output n115;
    output n7933;
    output n16276;
    output n80;
    output n16264;
    output n16336;
    output n7931;
    output n16265;
    output n117;
    output n16421;
    
    wire clk_in_c /* synthesis SET_AS_NETWORK=clk_in_c, is_clock=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(9[8:14])
    wire [17:0]instruction_c /* synthesis syn_ramstyle="block_ram", ram_style="distributed" */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    wire [17:0]n804;
    wire [17:0]n747;
    wire [17:0]n690;
    wire [17:0]n785;
    wire [17:0]n576;
    wire [17:0]n728;
    wire [17:0]n671;
    wire [17:0]n557;
    
    wire n19804, n19805, n19811, n19812, n19818, n19819, n19825, 
        n19826, n19832, n19833, n199, n236, n19839, n19840, n19922, 
        n19921, n19920, n19919, n19915, n19914, n19913, n19912, 
        n19908, n19907, n19846, n19847, n19906, n19905, n19901, 
        n19900, n19899, n19898, n19894, n19893, n19892, n19891, 
        n19887, n19886, n19885, n19884, n19880, n19879, n19878, 
        n19877, n19873, n19872, n19871, n19853, n19854, n19870, 
        n19866, n19865, n19864, n19863, n19859, n16465, n19858, 
        n19857, n19856, n19852, n19851, n19850, n19849, n19845, 
        n19844, n19843, n19842, n19838, n19837, n19860, n19861, 
        n19836, n19835, n19831, n19830, n210, n19829, n19828, 
        n19824, n19823, n19822, n19821, n19817, n19816, n19815, 
        n19814, n19867, n19868, n19810, n19809, n19808, n19807, 
        n19803, n19802, n19801, n19800, n19874, n19875, n19881, 
        n19882, n19888, n19889, n19916, n19917, n19895, n19896, 
        n19923, n19924, n19902, n19903, n19909, n19910;
    
    PDPW8KC mux_133 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
            .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), .DI11(GND_net), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(GND_net), .ADW1(GND_net), 
            .ADW2(GND_net), .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), 
            .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), 
            .BE1(GND_net), .CEW(VCC_net), .CLKW(GND_net), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(address[0]), .ADR5(address[1]), 
            .ADR6(address[2]), .ADR7(address[3]), .ADR8(address[4]), .ADR9(address[5]), 
            .ADR10(address[6]), .ADR11(address[7]), .ADR12(address[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(clk_in_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n804[9]), 
            .DO1(n804[10]), .DO2(n804[11]), .DO3(n804[12]), .DO4(n804[13]), 
            .DO5(n804[14]), .DO6(n804[15]), .DO7(n804[16]), .DO8(n804[17]), 
            .DO9(n804[0]), .DO10(n804[1]), .DO11(n804[2]), .DO12(n804[3]), 
            .DO13(n804[4]), .DO14(n804[5]), .DO15(n804[6]), .DO16(n804[7]), 
            .DO17(n804[8]));
    defparam mux_133.DATA_WIDTH_W = 18;
    defparam mux_133.DATA_WIDTH_R = 18;
    defparam mux_133.REGMODE = "NOREG";
    defparam mux_133.CSDECODE_W = "0b000";
    defparam mux_133.CSDECODE_R = "0b000";
    defparam mux_133.GSR = "DISABLED";
    defparam mux_133.RESETMODE = "ASYNC";
    defparam mux_133.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_133.INIT_DATA = "STATIC";
    defparam mux_133.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_133.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC mux_130 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
            .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), .DI11(GND_net), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(GND_net), .ADW1(GND_net), 
            .ADW2(GND_net), .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), 
            .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), 
            .BE1(GND_net), .CEW(VCC_net), .CLKW(GND_net), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(address[0]), .ADR5(address[1]), 
            .ADR6(address[2]), .ADR7(address[3]), .ADR8(address[4]), .ADR9(address[5]), 
            .ADR10(address[6]), .ADR11(address[7]), .ADR12(address[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(clk_in_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n747[9]), 
            .DO1(n747[10]), .DO2(n747[11]), .DO3(n747[12]), .DO4(n747[13]), 
            .DO5(n747[14]), .DO6(n747[15]), .DO7(n747[16]), .DO8(n747[17]), 
            .DO9(n747[0]), .DO10(n747[1]), .DO11(n747[2]), .DO12(n747[3]), 
            .DO13(n747[4]), .DO14(n747[5]), .DO15(n747[6]), .DO16(n747[7]), 
            .DO17(n747[8]));
    defparam mux_130.DATA_WIDTH_W = 18;
    defparam mux_130.DATA_WIDTH_R = 18;
    defparam mux_130.REGMODE = "NOREG";
    defparam mux_130.CSDECODE_W = "0b000";
    defparam mux_130.CSDECODE_R = "0b000";
    defparam mux_130.GSR = "DISABLED";
    defparam mux_130.RESETMODE = "ASYNC";
    defparam mux_130.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_130.INIT_DATA = "STATIC";
    defparam mux_130.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_130.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC mux_127 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
            .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), .DI11(GND_net), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(GND_net), .ADW1(GND_net), 
            .ADW2(GND_net), .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), 
            .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), 
            .BE1(GND_net), .CEW(VCC_net), .CLKW(GND_net), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(address[0]), .ADR5(address[1]), 
            .ADR6(address[2]), .ADR7(address[3]), .ADR8(address[4]), .ADR9(address[5]), 
            .ADR10(address[6]), .ADR11(address[7]), .ADR12(address[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(clk_in_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n690[9]), 
            .DO1(n690[10]), .DO2(n690[11]), .DO3(n690[12]), .DO4(n690[13]), 
            .DO5(n690[14]), .DO6(n690[15]), .DO7(n690[16]), .DO8(n690[17]), 
            .DO9(n690[0]), .DO10(n690[1]), .DO11(n690[2]), .DO12(n690[3]), 
            .DO13(n690[4]), .DO14(n690[5]), .DO15(n690[6]), .DO16(n690[7]), 
            .DO17(n690[8]));
    defparam mux_127.DATA_WIDTH_W = 18;
    defparam mux_127.DATA_WIDTH_R = 18;
    defparam mux_127.REGMODE = "NOREG";
    defparam mux_127.CSDECODE_W = "0b000";
    defparam mux_127.CSDECODE_R = "0b000";
    defparam mux_127.GSR = "DISABLED";
    defparam mux_127.RESETMODE = "ASYNC";
    defparam mux_127.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_127.INIT_DATA = "STATIC";
    defparam mux_127.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_127.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC mux_132 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
            .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), .DI11(GND_net), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(GND_net), .ADW1(GND_net), 
            .ADW2(GND_net), .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), 
            .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), 
            .BE1(GND_net), .CEW(VCC_net), .CLKW(GND_net), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(address[0]), .ADR5(address[1]), 
            .ADR6(address[2]), .ADR7(address[3]), .ADR8(address[4]), .ADR9(address[5]), 
            .ADR10(address[6]), .ADR11(address[7]), .ADR12(address[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(clk_in_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n785[9]), 
            .DO1(n785[10]), .DO2(n785[11]), .DO3(n785[12]), .DO4(n785[13]), 
            .DO5(n785[14]), .DO6(n785[15]), .DO7(n785[16]), .DO8(n785[17]), 
            .DO9(n785[0]), .DO10(n785[1]), .DO11(n785[2]), .DO12(n785[3]), 
            .DO13(n785[4]), .DO14(n785[5]), .DO15(n785[6]), .DO16(n785[7]), 
            .DO17(n785[8]));
    defparam mux_132.DATA_WIDTH_W = 18;
    defparam mux_132.DATA_WIDTH_R = 18;
    defparam mux_132.REGMODE = "NOREG";
    defparam mux_132.CSDECODE_W = "0b000";
    defparam mux_132.CSDECODE_R = "0b000";
    defparam mux_132.GSR = "DISABLED";
    defparam mux_132.RESETMODE = "ASYNC";
    defparam mux_132.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_132.INIT_DATA = "STATIC";
    defparam mux_132.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_132.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC mux_121 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
            .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), .DI11(GND_net), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(GND_net), .ADW1(GND_net), 
            .ADW2(GND_net), .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), 
            .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), 
            .BE1(GND_net), .CEW(VCC_net), .CLKW(GND_net), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(address[0]), .ADR5(address[1]), 
            .ADR6(address[2]), .ADR7(address[3]), .ADR8(address[4]), .ADR9(address[5]), 
            .ADR10(address[6]), .ADR11(address[7]), .ADR12(address[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(clk_in_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n576[9]), 
            .DO1(n576[10]), .DO2(n576[11]), .DO3(n576[12]), .DO4(n576[13]), 
            .DO5(n576[14]), .DO6(n576[15]), .DO7(n576[16]), .DO8(n576[17]), 
            .DO9(n576[0]), .DO10(n576[1]), .DO11(n576[2]), .DO12(n576[3]), 
            .DO13(n576[4]), .DO14(n576[5]), .DO15(n576[6]), .DO16(n576[7]), 
            .DO17(n576[8]));
    defparam mux_121.DATA_WIDTH_W = 18;
    defparam mux_121.DATA_WIDTH_R = 18;
    defparam mux_121.REGMODE = "NOREG";
    defparam mux_121.CSDECODE_W = "0b000";
    defparam mux_121.CSDECODE_R = "0b000";
    defparam mux_121.GSR = "DISABLED";
    defparam mux_121.RESETMODE = "ASYNC";
    defparam mux_121.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_121.INIT_DATA = "STATIC";
    defparam mux_121.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_121.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC mux_129 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
            .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), .DI11(GND_net), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(GND_net), .ADW1(GND_net), 
            .ADW2(GND_net), .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), 
            .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), 
            .BE1(GND_net), .CEW(VCC_net), .CLKW(GND_net), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(address[0]), .ADR5(address[1]), 
            .ADR6(address[2]), .ADR7(address[3]), .ADR8(address[4]), .ADR9(address[5]), 
            .ADR10(address[6]), .ADR11(address[7]), .ADR12(address[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(clk_in_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n728[9]), 
            .DO1(n728[10]), .DO2(n728[11]), .DO3(n728[12]), .DO4(n728[13]), 
            .DO5(n728[14]), .DO6(n728[15]), .DO7(n728[16]), .DO8(n728[17]), 
            .DO9(n728[0]), .DO10(n728[1]), .DO11(n728[2]), .DO12(n728[3]), 
            .DO13(n728[4]), .DO14(n728[5]), .DO15(n728[6]), .DO16(n728[7]), 
            .DO17(n728[8]));
    defparam mux_129.DATA_WIDTH_W = 18;
    defparam mux_129.DATA_WIDTH_R = 18;
    defparam mux_129.REGMODE = "NOREG";
    defparam mux_129.CSDECODE_W = "0b000";
    defparam mux_129.CSDECODE_R = "0b000";
    defparam mux_129.GSR = "DISABLED";
    defparam mux_129.RESETMODE = "ASYNC";
    defparam mux_129.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_129.INIT_DATA = "STATIC";
    defparam mux_129.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_129.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC mux_126 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
            .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), .DI11(GND_net), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(GND_net), .ADW1(GND_net), 
            .ADW2(GND_net), .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), 
            .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), 
            .BE1(GND_net), .CEW(VCC_net), .CLKW(GND_net), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(address[0]), .ADR5(address[1]), 
            .ADR6(address[2]), .ADR7(address[3]), .ADR8(address[4]), .ADR9(address[5]), 
            .ADR10(address[6]), .ADR11(address[7]), .ADR12(address[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(clk_in_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n671[9]), 
            .DO1(n671[10]), .DO2(n671[11]), .DO3(n671[12]), .DO4(n671[13]), 
            .DO5(n671[14]), .DO6(n671[15]), .DO7(n671[16]), .DO8(n671[17]), 
            .DO9(n671[0]), .DO10(n671[1]), .DO11(n671[2]), .DO12(n671[3]), 
            .DO13(n671[4]), .DO14(n671[5]), .DO15(n671[6]), .DO16(n671[7]), 
            .DO17(n671[8]));
    defparam mux_126.DATA_WIDTH_W = 18;
    defparam mux_126.DATA_WIDTH_R = 18;
    defparam mux_126.REGMODE = "NOREG";
    defparam mux_126.CSDECODE_W = "0b000";
    defparam mux_126.CSDECODE_R = "0b000";
    defparam mux_126.GSR = "DISABLED";
    defparam mux_126.RESETMODE = "ASYNC";
    defparam mux_126.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_126.INIT_DATA = "STATIC";
    defparam mux_126.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_126.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC mux_120 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
            .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), .DI11(GND_net), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(GND_net), .ADW1(GND_net), 
            .ADW2(GND_net), .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), 
            .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), 
            .BE1(GND_net), .CEW(VCC_net), .CLKW(GND_net), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(address[0]), .ADR5(address[1]), 
            .ADR6(address[2]), .ADR7(address[3]), .ADR8(address[4]), .ADR9(address[5]), 
            .ADR10(address[6]), .ADR11(address[7]), .ADR12(address[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(clk_in_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n557[9]), 
            .DO1(n557[10]), .DO2(n557[11]), .DO3(n557[12]), .DO4(n557[13]), 
            .DO5(n557[14]), .DO6(n557[15]), .DO7(n557[16]), .DO8(n557[17]), 
            .DO9(n557[0]), .DO10(n557[1]), .DO11(n557[2]), .DO12(n557[3]), 
            .DO13(n557[4]), .DO14(n557[5]), .DO15(n557[6]), .DO16(n557[7]), 
            .DO17(n557[8]));
    defparam mux_120.DATA_WIDTH_W = 18;
    defparam mux_120.DATA_WIDTH_R = 18;
    defparam mux_120.REGMODE = "NOREG";
    defparam mux_120.CSDECODE_W = "0b000";
    defparam mux_120.CSDECODE_R = "0b000";
    defparam mux_120.GSR = "DISABLED";
    defparam mux_120.RESETMODE = "ASYNC";
    defparam mux_120.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_120.INIT_DATA = "STATIC";
    defparam mux_120.INITVAL_00 = "0x14D063E02214D063E02914D0609D002800109D002DC0201C072DB002FB0001B662FA012DA0101AFE";
    defparam mux_120.INITVAL_01 = "0x01E013A00A0DE2009E00200302200A2FE0001E003A00A0DE1009E00200302200A3E01414D063E01B";
    defparam mux_120.INITVAL_02 = "0x2200A2FE0001E033A00A0DE8009E00200302200A2FE0001E023A00A0DE4009E00200302200A2FE00";
    defparam mux_120.INITVAL_03 = "0x11C010BC0025000360381B2001B10019001000002203801080011A90120322038010E00112E01200";
    defparam mux_120.INITVAL_04 = "0x2DA0114A0C0BA01250002FC002DC0001C003604A1DBA003BF000BC011C063604A1DB0A03B0F00BC0";
    defparam mux_120.INITVAL_05 = "0x0000000000000000000000000000000000000000290012003E2004D280000000000000250002FA01";
    defparam mux_120.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_120.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    L6MUX21 i16636 (.D0(n19804), .D1(n19805), .SD(address[11]), .Z(instruction[0]));
    L6MUX21 i16643 (.D0(n19811), .D1(n19812), .SD(address[11]), .Z(instruction[1]));
    L6MUX21 i16650 (.D0(n19818), .D1(n19819), .SD(address[11]), .Z(instruction[2]));
    L6MUX21 i16657 (.D0(n19825), .D1(n19826), .SD(address[11]), .Z(instruction[3]));
    L6MUX21 i16664 (.D0(n19832), .D1(n19833), .SD(address[11]), .Z(instruction[4]));
    LUT4 i1_2_lut_3_lut_4_lut (.A(n199), .B(n236), .C(n16312), .D(n11778), 
         .Z(n16351)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_204 (.A(n199), .B(n236), .C(n11714), 
         .D(n11778), .Z(n16261)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_204.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_adj_205 (.A(n199), .B(n236), .C(n7908), 
         .D(n16392), .Z(n7941)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_205.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_206 (.A(n199), .B(n236), .C(n7762), 
         .D(n7726), .Z(n82)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_206.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_207 (.A(n199), .B(n236), .C(n7762), 
         .D(n16392), .Z(n81)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_207.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_208 (.A(n199), .B(n236), .C(n16312), 
         .D(n7876), .Z(n16315)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_208.init = 16'h2000;
    L6MUX21 i16671 (.D0(n19839), .D1(n19840), .SD(address[11]), .Z(instruction[5]));
    LUT4 i1_2_lut_rep_542_4_lut (.A(instruction[0]), .B(n16417), .C(instruction[2]), 
         .D(instruction[1]), .Z(n22109)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_542_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_3_lut (.A(instruction[0]), .B(n7646), .C(instruction[3]), 
         .Z(n199)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h0404;
    LUT4 i1_3_lut_3_lut (.A(instruction[2]), .B(instruction[1]), .C(n199), 
         .Z(n2075)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_209 (.A(n199), .B(instruction[1]), .C(instruction[2]), 
         .D(n7876), .Z(n9)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_209.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_210 (.A(n199), .B(instruction[1]), .C(instruction[2]), 
         .D(n7726), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_210.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_211 (.A(n199), .B(instruction[1]), .C(instruction[2]), 
         .D(n11778), .Z(n8)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_211.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_212 (.A(n199), .B(instruction[1]), .C(instruction[2]), 
         .D(n16392), .Z(n7)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_212.init = 16'h8000;
    LUT4 i16752_3_lut (.A(n785[17]), .B(n804[17]), .C(address[9]), .Z(n19922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16752_3_lut.init = 16'hcaca;
    LUT4 i16751_3_lut (.A(n671[17]), .B(n690[17]), .C(address[9]), .Z(n19921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16751_3_lut.init = 16'hcaca;
    LUT4 i16750_3_lut (.A(n728[17]), .B(n747[17]), .C(address[9]), .Z(n19920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16750_3_lut.init = 16'hcaca;
    LUT4 i16749_3_lut (.A(n557[17]), .B(n576[17]), .C(address[9]), .Z(n19919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16749_3_lut.init = 16'hcaca;
    LUT4 i16745_3_lut (.A(n785[16]), .B(n804[16]), .C(address[9]), .Z(n19915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16745_3_lut.init = 16'hcaca;
    LUT4 i16744_3_lut (.A(n671[16]), .B(n690[16]), .C(address[9]), .Z(n19914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16744_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_213 (.A(n199), .B(n236), .C(n7762), 
         .D(n11778), .Z(n83)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_213.init = 16'h0020;
    LUT4 i16743_3_lut (.A(n728[16]), .B(n747[16]), .C(address[9]), .Z(n19913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16743_3_lut.init = 16'hcaca;
    LUT4 i16742_3_lut (.A(n557[16]), .B(n576[16]), .C(address[9]), .Z(n19912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16742_3_lut.init = 16'hcaca;
    LUT4 i16738_3_lut (.A(n785[15]), .B(n804[15]), .C(address[9]), .Z(n19908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16738_3_lut.init = 16'hcaca;
    LUT4 i16737_3_lut (.A(n671[15]), .B(n690[15]), .C(address[9]), .Z(n19907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16737_3_lut.init = 16'hcaca;
    L6MUX21 i16678 (.D0(n19846), .D1(n19847), .SD(address[11]), .Z(instruction[6]));
    LUT4 i16736_3_lut (.A(n728[15]), .B(n747[15]), .C(address[9]), .Z(n19906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16736_3_lut.init = 16'hcaca;
    LUT4 i16735_3_lut (.A(n557[15]), .B(n576[15]), .C(address[9]), .Z(n19905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16735_3_lut.init = 16'hcaca;
    LUT4 i16731_3_lut (.A(n785[14]), .B(n804[14]), .C(address[9]), .Z(n19901)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16731_3_lut.init = 16'hcaca;
    LUT4 i16730_3_lut (.A(n671[14]), .B(n690[14]), .C(address[9]), .Z(n19900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16730_3_lut.init = 16'hcaca;
    LUT4 i16729_3_lut (.A(n728[14]), .B(n747[14]), .C(address[9]), .Z(n19899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16729_3_lut.init = 16'hcaca;
    LUT4 i16728_3_lut (.A(n557[14]), .B(n576[14]), .C(address[9]), .Z(n19898)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16728_3_lut.init = 16'hcaca;
    LUT4 i16724_3_lut (.A(n785[13]), .B(n804[13]), .C(address[9]), .Z(n19894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16724_3_lut.init = 16'hcaca;
    LUT4 i16723_3_lut (.A(n671[13]), .B(n690[13]), .C(address[9]), .Z(n19893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16723_3_lut.init = 16'hcaca;
    LUT4 i16722_3_lut (.A(n728[13]), .B(n747[13]), .C(address[9]), .Z(n19892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16722_3_lut.init = 16'hcaca;
    LUT4 i16721_3_lut (.A(n557[13]), .B(n576[13]), .C(address[9]), .Z(n19891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16721_3_lut.init = 16'hcaca;
    LUT4 i16717_3_lut (.A(n785[12]), .B(n804[12]), .C(address[9]), .Z(n19887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16717_3_lut.init = 16'hcaca;
    LUT4 i16716_3_lut (.A(n671[12]), .B(n690[12]), .C(address[9]), .Z(n19886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16716_3_lut.init = 16'hcaca;
    LUT4 i16715_3_lut (.A(n728[12]), .B(n747[12]), .C(address[9]), .Z(n19885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16715_3_lut.init = 16'hcaca;
    LUT4 i16714_3_lut (.A(n557[12]), .B(n576[12]), .C(address[9]), .Z(n19884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16714_3_lut.init = 16'hcaca;
    LUT4 i16710_3_lut (.A(n785[11]), .B(n804[11]), .C(address[9]), .Z(n19880)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16710_3_lut.init = 16'hcaca;
    LUT4 i16709_3_lut (.A(n671[11]), .B(n690[11]), .C(address[9]), .Z(n19879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16709_3_lut.init = 16'hcaca;
    LUT4 i16708_3_lut (.A(n728[11]), .B(n747[11]), .C(address[9]), .Z(n19878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16708_3_lut.init = 16'hcaca;
    LUT4 i16707_3_lut (.A(n557[11]), .B(n576[11]), .C(address[9]), .Z(n19877)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16707_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_214 (.A(n199), .B(n236), .C(n7908), 
         .D(n7726), .Z(n7940)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_214.init = 16'h2000;
    LUT4 i16703_3_lut (.A(n785[10]), .B(n804[10]), .C(address[9]), .Z(n19873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16703_3_lut.init = 16'hcaca;
    LUT4 i16702_3_lut (.A(n671[10]), .B(n690[10]), .C(address[9]), .Z(n19872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16702_3_lut.init = 16'hcaca;
    LUT4 i16701_3_lut (.A(n728[10]), .B(n747[10]), .C(address[9]), .Z(n19871)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16701_3_lut.init = 16'hcaca;
    L6MUX21 i16685 (.D0(n19853), .D1(n19854), .SD(address[11]), .Z(instruction[7]));
    LUT4 i1_2_lut_3_lut_4_lut_adj_215 (.A(n199), .B(n236), .C(n7908), 
         .D(n7876), .Z(n7942)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_215.init = 16'h2000;
    LUT4 i16700_3_lut (.A(n557[10]), .B(n576[10]), .C(address[9]), .Z(n19870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16700_3_lut.init = 16'hcaca;
    LUT4 i16696_3_lut (.A(n785[9]), .B(n804[9]), .C(address[9]), .Z(n19866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16696_3_lut.init = 16'hcaca;
    LUT4 i16695_3_lut (.A(n671[9]), .B(n690[9]), .C(address[9]), .Z(n19865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16695_3_lut.init = 16'hcaca;
    LUT4 i16694_3_lut (.A(n728[9]), .B(n747[9]), .C(address[9]), .Z(n19864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16694_3_lut.init = 16'hcaca;
    LUT4 i16693_3_lut (.A(n557[9]), .B(n576[9]), .C(address[9]), .Z(n19863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16693_3_lut.init = 16'hcaca;
    LUT4 i16689_3_lut (.A(n785[8]), .B(n804[8]), .C(address[9]), .Z(n19859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16689_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_216 (.A(instruction[0]), .B(instruction[1]), 
         .C(instruction[2]), .Z(n16465)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_216.init = 16'h8080;
    LUT4 i2_3_lut_4_lut (.A(instruction[2]), .B(instruction[0]), .C(n16417), 
         .D(instruction[1]), .Z(n2081)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h1000;
    LUT4 i16688_3_lut (.A(n671[8]), .B(n690[8]), .C(address[9]), .Z(n19858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16688_3_lut.init = 16'hcaca;
    LUT4 i16687_3_lut (.A(n728[8]), .B(n747[8]), .C(address[9]), .Z(n19857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16687_3_lut.init = 16'hcaca;
    LUT4 i16686_3_lut (.A(n557[8]), .B(n576[8]), .C(address[9]), .Z(n19856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16686_3_lut.init = 16'hcaca;
    LUT4 i16682_3_lut (.A(n785[7]), .B(n804[7]), .C(address[9]), .Z(n19852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16682_3_lut.init = 16'hcaca;
    LUT4 i16681_3_lut (.A(n671[7]), .B(n690[7]), .C(address[9]), .Z(n19851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16681_3_lut.init = 16'hcaca;
    LUT4 i16680_3_lut (.A(n728[7]), .B(n747[7]), .C(address[9]), .Z(n19850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16680_3_lut.init = 16'hcaca;
    LUT4 i16679_3_lut (.A(n557[7]), .B(n576[7]), .C(address[9]), .Z(n19849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16679_3_lut.init = 16'hcaca;
    LUT4 i16675_3_lut (.A(n785[6]), .B(n804[6]), .C(address[9]), .Z(n19845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16675_3_lut.init = 16'hcaca;
    LUT4 i16674_3_lut (.A(n671[6]), .B(n690[6]), .C(address[9]), .Z(n19844)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16674_3_lut.init = 16'hcaca;
    LUT4 i16673_3_lut (.A(n728[6]), .B(n747[6]), .C(address[9]), .Z(n19843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16673_3_lut.init = 16'hcaca;
    LUT4 i16672_3_lut (.A(n557[6]), .B(n576[6]), .C(address[9]), .Z(n19842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16672_3_lut.init = 16'hcaca;
    LUT4 i16668_3_lut (.A(n785[5]), .B(n804[5]), .C(address[9]), .Z(n19838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16668_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_217 (.A(n199), .B(n236), .C(n16312), 
         .D(n16392), .Z(n16348)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_217.init = 16'h2000;
    LUT4 i16667_3_lut (.A(n671[5]), .B(n690[5]), .C(address[9]), .Z(n19837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16667_3_lut.init = 16'hcaca;
    L6MUX21 i16692 (.D0(n19860), .D1(n19861), .SD(address[11]), .Z(instruction[8]));
    LUT4 i16666_3_lut (.A(n728[5]), .B(n747[5]), .C(address[9]), .Z(n19836)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16666_3_lut.init = 16'hcaca;
    LUT4 i16665_3_lut (.A(n557[5]), .B(n576[5]), .C(address[9]), .Z(n19835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16665_3_lut.init = 16'hcaca;
    LUT4 i16661_3_lut (.A(n785[4]), .B(n804[4]), .C(address[9]), .Z(n19831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16661_3_lut.init = 16'hcaca;
    LUT4 i16660_3_lut (.A(n671[4]), .B(n690[4]), .C(address[9]), .Z(n19830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16660_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_218 (.A(instruction[0]), .B(instruction[3]), 
         .C(n7646), .Z(n210)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_218.init = 16'h4040;
    LUT4 i16659_3_lut (.A(n728[4]), .B(n747[4]), .C(address[9]), .Z(n19829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16659_3_lut.init = 16'hcaca;
    LUT4 i16658_3_lut (.A(n557[4]), .B(n576[4]), .C(address[9]), .Z(n19828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16658_3_lut.init = 16'hcaca;
    LUT4 i16654_3_lut (.A(n785[3]), .B(n804[3]), .C(address[9]), .Z(n19824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16654_3_lut.init = 16'hcaca;
    LUT4 i16653_3_lut (.A(n671[3]), .B(n690[3]), .C(address[9]), .Z(n19823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16653_3_lut.init = 16'hcaca;
    LUT4 i16652_3_lut (.A(n728[3]), .B(n747[3]), .C(address[9]), .Z(n19822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16652_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_219 (.A(n7646), .B(instruction[3]), .C(n16465), 
         .D(n7876), .Z(n9_adj_6)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_219.init = 16'h2000;
    LUT4 i16651_3_lut (.A(n557[3]), .B(n576[3]), .C(address[9]), .Z(n19821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16651_3_lut.init = 16'hcaca;
    LUT4 i16647_3_lut (.A(n785[2]), .B(n804[2]), .C(address[9]), .Z(n19817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16647_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_220 (.A(n7646), .B(instruction[3]), .C(n16465), 
         .D(n7726), .Z(n10_adj_7)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_220.init = 16'h2000;
    LUT4 i16646_3_lut (.A(n671[2]), .B(n690[2]), .C(address[9]), .Z(n19816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16646_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_221 (.A(n7646), .B(instruction[3]), .C(n16465), 
         .D(n16392), .Z(n7_adj_8)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_221.init = 16'h2000;
    LUT4 i16645_3_lut (.A(n728[2]), .B(n747[2]), .C(address[9]), .Z(n19815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16645_3_lut.init = 16'hcaca;
    LUT4 i16644_3_lut (.A(n557[2]), .B(n576[2]), .C(address[9]), .Z(n19814)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16644_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_222 (.A(n7646), .B(instruction[3]), .C(n16465), 
         .D(n11778), .Z(n8_adj_9)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_222.init = 16'h0020;
    L6MUX21 i16699 (.D0(n19867), .D1(n19868), .SD(address[11]), .Z(instruction[9]));
    LUT4 i16640_3_lut (.A(n785[1]), .B(n804[1]), .C(address[9]), .Z(n19810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16640_3_lut.init = 16'hcaca;
    LUT4 i16639_3_lut (.A(n671[1]), .B(n690[1]), .C(address[9]), .Z(n19809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16639_3_lut.init = 16'hcaca;
    LUT4 i16638_3_lut (.A(n728[1]), .B(n747[1]), .C(address[9]), .Z(n19808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16638_3_lut.init = 16'hcaca;
    LUT4 i16637_3_lut (.A(n557[1]), .B(n576[1]), .C(address[9]), .Z(n19807)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16637_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_223 (.A(n199), .B(n236), .C(n11714), 
         .D(n7726), .Z(n16277)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_223.init = 16'h0200;
    LUT4 i16633_3_lut (.A(n785[0]), .B(n804[0]), .C(address[9]), .Z(n19803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16633_3_lut.init = 16'hcaca;
    LUT4 i16632_3_lut (.A(n671[0]), .B(n690[0]), .C(address[9]), .Z(n19802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16632_3_lut.init = 16'hcaca;
    LUT4 i16631_3_lut (.A(n728[0]), .B(n747[0]), .C(address[9]), .Z(n19801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16631_3_lut.init = 16'hcaca;
    LUT4 i16630_3_lut (.A(n557[0]), .B(n576[0]), .C(address[9]), .Z(n19800)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16630_3_lut.init = 16'hcaca;
    L6MUX21 i16706 (.D0(n19874), .D1(n19875), .SD(address[11]), .Z(instruction[10]));
    L6MUX21 i16713 (.D0(n19881), .D1(n19882), .SD(address[11]), .Z(instruction[11]));
    LUT4 i1_2_lut_3_lut_4_lut_adj_224 (.A(n199), .B(n236), .C(n7908), 
         .D(n11778), .Z(n7939)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_224.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_225 (.A(n16417), .B(n16465), .C(n11714), 
         .D(n7726), .Z(n16289)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_225.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_226 (.A(n16417), .B(n16465), .C(n7908), 
         .D(n7726), .Z(n7921)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_226.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_227 (.A(n16417), .B(n16465), .C(n16312), 
         .D(n7876), .Z(n16345)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_227.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_228 (.A(n16417), .B(n16465), .C(n7908), 
         .D(n7876), .Z(n7919)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_228.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_229 (.A(n16417), .B(n16465), .C(n11714), 
         .D(n16392), .Z(n16285)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_229.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_230 (.A(n16417), .B(n16465), .C(n16312), 
         .D(n16392), .Z(n16332)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_230.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_231 (.A(n16417), .B(n16465), .C(n7762), 
         .D(n7726), .Z(n145)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_231.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_232 (.A(n16417), .B(n16465), .C(n11714), 
         .D(n11778), .Z(n16284)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_232.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_233 (.A(n16417), .B(n16465), .C(n16312), 
         .D(n11778), .Z(n16327)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_233.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_234 (.A(n16417), .B(n16465), .C(n7908), 
         .D(n16392), .Z(n7920)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_234.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_235 (.A(n16417), .B(n16465), .C(n7762), 
         .D(n16392), .Z(n143)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_235.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_236 (.A(n16417), .B(n16465), .C(n7762), 
         .D(n7876), .Z(n142)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_236.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_237 (.A(n16417), .B(n16465), .C(n11714), 
         .D(n7876), .Z(n16290)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_237.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_238 (.A(n16417), .B(n16465), .C(n16312), 
         .D(n7726), .Z(n16346)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_238.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_239 (.A(n16417), .B(n16465), .C(n7908), 
         .D(n11778), .Z(n7922)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_239.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_240 (.A(n16417), .B(n16465), .C(n7762), 
         .D(n11778), .Z(n146)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_240.init = 16'h0080;
    L6MUX21 i16720 (.D0(n19888), .D1(n19889), .SD(address[11]), .Z(instruction[12]));
    LUT4 i1_3_lut (.A(instruction[2]), .B(instruction[1]), .C(n199), .Z(n2071)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_241 (.A(n210), .B(instruction[2]), .C(instruction[1]), 
         .D(n11778), .Z(n8_adj_10)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_241.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_adj_242 (.A(n199), .B(n236), .C(n16312), 
         .D(n7726), .Z(n16316)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_242.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_243 (.A(n199), .B(n236), .C(n11714), 
         .D(n16392), .Z(n16260)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_243.init = 16'h0200;
    LUT4 i2_3_lut (.A(instruction[2]), .B(n210), .C(instruction[1]), .Z(n2085)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i2_3_lut.init = 16'h0808;
    LUT4 i1_2_lut (.A(instruction[3]), .B(n7646), .Z(n16417)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_244 (.A(n206), .B(n210), .C(n7762), 
         .D(n7726), .Z(n116)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_244.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_245 (.A(n206), .B(n210), .C(n16312), 
         .D(n7726), .Z(n16319)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_245.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_246 (.A(n206), .B(n210), .C(n7908), 
         .D(n7876), .Z(n7934)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_246.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_247 (.A(n206), .B(n210), .C(n11714), 
         .D(n7726), .Z(n16279)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_247.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_248 (.A(n206), .B(n210), .C(n7908), 
         .D(n7726), .Z(n7932)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_248.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_249 (.A(n206), .B(n210), .C(n7762), 
         .D(n7876), .Z(n114)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_249.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_250 (.A(n206), .B(n210), .C(n16312), 
         .D(n7876), .Z(n16318)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_250.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_251 (.A(n206), .B(n210), .C(n11714), 
         .D(n7876), .Z(n16278)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_251.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_252 (.A(n206), .B(n210), .C(n16312), 
         .D(n16392), .Z(n16330)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_252.init = 16'h8000;
    L6MUX21 i16748 (.D0(n19916), .D1(n19917), .SD(address[11]), .Z(instruction[16]));
    LUT4 i1_2_lut_3_lut_4_lut_adj_253 (.A(n206), .B(n210), .C(n7762), 
         .D(n16392), .Z(n115)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_253.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_254 (.A(n206), .B(n210), .C(n7908), 
         .D(n16392), .Z(n7933)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_254.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_255 (.A(n199), .B(n236), .C(n11714), 
         .D(n7876), .Z(n16276)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_255.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_256 (.A(n199), .B(n236), .C(n7762), 
         .D(n7876), .Z(n80)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_256.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_257 (.A(n206), .B(n210), .C(n11714), 
         .D(n16392), .Z(n16264)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_257.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_258 (.A(n206), .B(n210), .C(n16312), 
         .D(n11778), .Z(n16336)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_258.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_259 (.A(n206), .B(n210), .C(n7908), 
         .D(n11778), .Z(n7931)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_259.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_260 (.A(n206), .B(n210), .C(n11714), 
         .D(n11778), .Z(n16265)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_260.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_261 (.A(n206), .B(n210), .C(n7762), 
         .D(n11778), .Z(n117)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_261.init = 16'h0080;
    L6MUX21 i16727 (.D0(n19895), .D1(n19896), .SD(address[11]), .Z(instruction[13]));
    L6MUX21 i16755 (.D0(n19923), .D1(n19924), .SD(address[11]), .Z(instruction[17]));
    LUT4 i1_2_lut_adj_262 (.A(n7646), .B(instruction[3]), .Z(n16421)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_262.init = 16'h2222;
    LUT4 i225_2_lut (.A(instruction[2]), .B(instruction[1]), .Z(n236)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i225_2_lut.init = 16'heeee;
    L6MUX21 i16734 (.D0(n19902), .D1(n19903), .SD(address[11]), .Z(instruction[14]));
    PFUMX i16634 (.BLUT(n19800), .ALUT(n19801), .C0(address[10]), .Z(n19804));
    PFUMX i16635 (.BLUT(n19802), .ALUT(n19803), .C0(address[10]), .Z(n19805));
    PFUMX i16641 (.BLUT(n19807), .ALUT(n19808), .C0(address[10]), .Z(n19811));
    PFUMX i16642 (.BLUT(n19809), .ALUT(n19810), .C0(address[10]), .Z(n19812));
    PFUMX i16648 (.BLUT(n19814), .ALUT(n19815), .C0(address[10]), .Z(n19818));
    PFUMX i16649 (.BLUT(n19816), .ALUT(n19817), .C0(address[10]), .Z(n19819));
    PFUMX i16655 (.BLUT(n19821), .ALUT(n19822), .C0(address[10]), .Z(n19825));
    PFUMX i16656 (.BLUT(n19823), .ALUT(n19824), .C0(address[10]), .Z(n19826));
    PFUMX i16662 (.BLUT(n19828), .ALUT(n19829), .C0(address[10]), .Z(n19832));
    PFUMX i16663 (.BLUT(n19830), .ALUT(n19831), .C0(address[10]), .Z(n19833));
    PFUMX i16669 (.BLUT(n19835), .ALUT(n19836), .C0(address[10]), .Z(n19839));
    PFUMX i16670 (.BLUT(n19837), .ALUT(n19838), .C0(address[10]), .Z(n19840));
    PFUMX i16676 (.BLUT(n19842), .ALUT(n19843), .C0(address[10]), .Z(n19846));
    PFUMX i16677 (.BLUT(n19844), .ALUT(n19845), .C0(address[10]), .Z(n19847));
    PFUMX i16683 (.BLUT(n19849), .ALUT(n19850), .C0(address[10]), .Z(n19853));
    PFUMX i16684 (.BLUT(n19851), .ALUT(n19852), .C0(address[10]), .Z(n19854));
    PFUMX i16690 (.BLUT(n19856), .ALUT(n19857), .C0(address[10]), .Z(n19860));
    PFUMX i16691 (.BLUT(n19858), .ALUT(n19859), .C0(address[10]), .Z(n19861));
    PFUMX i16697 (.BLUT(n19863), .ALUT(n19864), .C0(address[10]), .Z(n19867));
    PFUMX i16698 (.BLUT(n19865), .ALUT(n19866), .C0(address[10]), .Z(n19868));
    PFUMX i16704 (.BLUT(n19870), .ALUT(n19871), .C0(address[10]), .Z(n19874));
    PFUMX i16705 (.BLUT(n19872), .ALUT(n19873), .C0(address[10]), .Z(n19875));
    PFUMX i16711 (.BLUT(n19877), .ALUT(n19878), .C0(address[10]), .Z(n19881));
    PFUMX i16712 (.BLUT(n19879), .ALUT(n19880), .C0(address[10]), .Z(n19882));
    L6MUX21 i16741 (.D0(n19909), .D1(n19910), .SD(address[11]), .Z(instruction[15]));
    PFUMX i16718 (.BLUT(n19884), .ALUT(n19885), .C0(address[10]), .Z(n19888));
    PFUMX i16719 (.BLUT(n19886), .ALUT(n19887), .C0(address[10]), .Z(n19889));
    PFUMX i16725 (.BLUT(n19891), .ALUT(n19892), .C0(address[10]), .Z(n19895));
    PFUMX i16726 (.BLUT(n19893), .ALUT(n19894), .C0(address[10]), .Z(n19896));
    PFUMX i16732 (.BLUT(n19898), .ALUT(n19899), .C0(address[10]), .Z(n19902));
    PFUMX i16733 (.BLUT(n19900), .ALUT(n19901), .C0(address[10]), .Z(n19903));
    PFUMX i16739 (.BLUT(n19905), .ALUT(n19906), .C0(address[10]), .Z(n19909));
    PFUMX i16740 (.BLUT(n19907), .ALUT(n19908), .C0(address[10]), .Z(n19910));
    PFUMX i16746 (.BLUT(n19912), .ALUT(n19913), .C0(address[10]), .Z(n19916));
    PFUMX i16747 (.BLUT(n19914), .ALUT(n19915), .C0(address[10]), .Z(n19917));
    PFUMX i16753 (.BLUT(n19919), .ALUT(n19920), .C0(address[10]), .Z(n19923));
    PFUMX i16754 (.BLUT(n19921), .ALUT(n19922), .C0(address[10]), .Z(n19924));
    
endmodule
//
// Verilog Description of module seg_display
//

module seg_display (seg_data_1, seg_led_1_c_5, seg_led_1_c_6, seg_led_1_c_1, 
            seg_led_1_c_2, seg_led_1_c_3, seg_data_2, seg_led_2_c_2, 
            seg_led_2_c_5, seg_led_2_c_6, seg_led_2_c_1, seg_led_2_c_3, 
            seg_led_2_c_0, seg_led_2_c_4, seg_led_1_c_0, seg_led_1_c_4) /* synthesis syn_module_defined=1 */ ;
    input [3:0]seg_data_1;
    output seg_led_1_c_5;
    output seg_led_1_c_6;
    output seg_led_1_c_1;
    output seg_led_1_c_2;
    output seg_led_1_c_3;
    input [3:0]seg_data_2;
    output seg_led_2_c_2;
    output seg_led_2_c_5;
    output seg_led_2_c_6;
    output seg_led_2_c_1;
    output seg_led_2_c_3;
    output seg_led_2_c_0;
    output seg_led_2_c_4;
    output seg_led_1_c_0;
    output seg_led_1_c_4;
    
    
    LUT4 seg_data_1_0__bdd_4_lut_18104 (.A(seg_data_1[0]), .B(seg_data_1[3]), 
         .C(seg_data_1[2]), .D(seg_data_1[1]), .Z(seg_led_1_c_5)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam seg_data_1_0__bdd_4_lut_18104.init = 16'h103d;
    LUT4 seg_data_1_1__bdd_4_lut (.A(seg_data_1[1]), .B(seg_data_1[3]), 
         .C(seg_data_1[0]), .D(seg_data_1[2]), .Z(seg_led_1_c_6)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B (D)+!B !(D)))) */ ;
    defparam seg_data_1_1__bdd_4_lut.init = 16'h1366;
    LUT4 seg_data_1_0__bdd_4_lut (.A(seg_data_1[0]), .B(seg_data_1[3]), 
         .C(seg_data_1[2]), .D(seg_data_1[1]), .Z(seg_led_1_c_1)) /* synthesis lut_function=(!(A (B (C+(D))+!B !((D)+!C))+!A (B (C+(D))+!B (C (D))))) */ ;
    defparam seg_data_1_0__bdd_4_lut.init = 16'h231f;
    LUT4 seg_data_1_2__bdd_4_lut (.A(seg_data_1[2]), .B(seg_data_1[0]), 
         .C(seg_data_1[3]), .D(seg_data_1[1]), .Z(seg_led_1_c_2)) /* synthesis lut_function=(!(A (C)+!A (B (C (D))+!B (D)))) */ ;
    defparam seg_data_1_2__bdd_4_lut.init = 16'h0e5f;
    LUT4 seg_data_1_3__bdd_4_lut (.A(seg_data_1[3]), .B(seg_data_1[0]), 
         .C(seg_data_1[2]), .D(seg_data_1[1]), .Z(seg_led_1_c_3)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam seg_data_1_3__bdd_4_lut.init = 16'h154b;
    LUT4 seg_data_2_2__bdd_4_lut (.A(seg_data_2[2]), .B(seg_data_2[0]), 
         .C(seg_data_2[3]), .D(seg_data_2[1]), .Z(seg_led_2_c_2)) /* synthesis lut_function=(!(A (C)+!A (B (C (D))+!B (D)))) */ ;
    defparam seg_data_2_2__bdd_4_lut.init = 16'h0e5f;
    LUT4 seg_data_2_0__bdd_4_lut_18112 (.A(seg_data_2[0]), .B(seg_data_2[3]), 
         .C(seg_data_2[2]), .D(seg_data_2[1]), .Z(seg_led_2_c_5)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam seg_data_2_0__bdd_4_lut_18112.init = 16'h103d;
    LUT4 seg_data_2_1__bdd_4_lut (.A(seg_data_2[1]), .B(seg_data_2[3]), 
         .C(seg_data_2[0]), .D(seg_data_2[2]), .Z(seg_led_2_c_6)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B (D)+!B !(D)))) */ ;
    defparam seg_data_2_1__bdd_4_lut.init = 16'h1366;
    LUT4 seg_data_2_0__bdd_4_lut (.A(seg_data_2[0]), .B(seg_data_2[3]), 
         .C(seg_data_2[2]), .D(seg_data_2[1]), .Z(seg_led_2_c_1)) /* synthesis lut_function=(!(A (B (C+(D))+!B !((D)+!C))+!A (B (C+(D))+!B (C (D))))) */ ;
    defparam seg_data_2_0__bdd_4_lut.init = 16'h231f;
    LUT4 seg_data_2_3__bdd_4_lut (.A(seg_data_2[3]), .B(seg_data_2[0]), 
         .C(seg_data_2[2]), .D(seg_data_2[1]), .Z(seg_led_2_c_3)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam seg_data_2_3__bdd_4_lut.init = 16'h154b;
    LUT4 mux_113_Mux_0_i15_4_lut (.A(seg_data_2[0]), .B(seg_data_2[2]), 
         .C(seg_data_2[3]), .D(seg_data_2[1]), .Z(seg_led_2_c_0)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/seg_display.v(30[28:43])
    defparam mux_113_Mux_0_i15_4_lut.init = 16'h0f39;
    LUT4 i17789_4_lut (.A(seg_data_2[0]), .B(seg_data_2[2]), .C(seg_data_2[3]), 
         .D(seg_data_2[1]), .Z(seg_led_2_c_4)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B (C (D))))) */ ;
    defparam i17789_4_lut.init = 16'h0511;
    LUT4 mux_112_Mux_0_i15_4_lut (.A(seg_data_1[0]), .B(seg_data_1[2]), 
         .C(seg_data_1[3]), .D(seg_data_1[1]), .Z(seg_led_1_c_0)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/seg_display.v(29[28:43])
    defparam mux_112_Mux_0_i15_4_lut.init = 16'h0f39;
    LUT4 i17786_4_lut (.A(seg_data_1[0]), .B(seg_data_1[2]), .C(seg_data_1[3]), 
         .D(seg_data_1[1]), .Z(seg_led_1_c_4)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B (C (D))))) */ ;
    defparam i17786_4_lut.init = 16'h0511;
    
endmodule
//
// Verilog Description of module mcu
//

module mcu (clk_in_c, n11714, instruction, n22301, interrupt, n16290, 
            out_port, port_id, write_strobe, GND_net, address, VCC_net, 
            n7762, n7908, n11778, n16278, n7876, n16417, n16279, 
            n206, n7646, n16312, n16392, n22109, n2085, n7921, 
            n2071, n2081, n7920, n7726, n7919, n16261, n16284, 
            n2075, n16277, n16260, n16285, n16276, n83, n146, 
            n16421, n82, n81, n143, n80, n16351, n16327, n16316, 
            n16348, n16332, rst_n_in, n16315, n7939, n7922, n7940, 
            n7941, n7942, n9, n9_adj_1, in_port, n7, n7_adj_2, 
            n10, n10_adj_3, n7931, n8, n8_adj_4, n16330, n16336, 
            n115, n117, n16264, n16265, n7934, n8_adj_5, n7933, 
            n7932, \cnt_p[22] , \cnt_p[23] , n14409, n857, n16289, 
            n16318, n16319, n114, n116, n145, n142, n16346, n16345) /* synthesis syn_module_defined=1 */ ;
    input clk_in_c;
    output n11714;
    input [17:0]instruction;
    output n22301;
    input interrupt;
    input n16290;
    output [7:0]out_port;
    output [7:0]port_id;
    output write_strobe;
    input GND_net;
    output [11:0]address;
    input VCC_net;
    output n7762;
    output n7908;
    output n11778;
    input n16278;
    output n7876;
    input n16417;
    input n16279;
    output n206;
    output n7646;
    output n16312;
    output n16392;
    input n22109;
    input n2085;
    input n7921;
    input n2071;
    input n2081;
    input n7920;
    output n7726;
    input n7919;
    input n16261;
    input n16284;
    input n2075;
    input n16277;
    input n16260;
    input n16285;
    input n16276;
    input n83;
    input n146;
    input n16421;
    input n82;
    input n81;
    input n143;
    input n80;
    input n16351;
    input n16327;
    input n16316;
    input n16348;
    input n16332;
    input rst_n_in;
    input n16315;
    input n7939;
    input n7922;
    input n7940;
    input n7941;
    input n7942;
    input n9;
    input n9_adj_1;
    input [7:0]in_port;
    input n7;
    input n7_adj_2;
    input n10;
    input n10_adj_3;
    input n7931;
    input n8;
    input n8_adj_4;
    input n16330;
    input n16336;
    input n115;
    input n117;
    input n16264;
    input n16265;
    input n7934;
    input n8_adj_5;
    input n7933;
    input n7932;
    input \cnt_p[22] ;
    input \cnt_p[23] ;
    input n14409;
    output n857;
    input n16289;
    input n16318;
    input n16319;
    input n114;
    input n116;
    input n145;
    input n142;
    input n16346;
    input n16345;
    
    wire clk_in_c /* synthesis SET_AS_NETWORK=clk_in_c, is_clock=1 */ ;   // f:/home/mini-mcu/step_fpga/top.v(9[8:14])
    wire [17:0]instruction_c /* synthesis syn_ramstyle="block_ram", ram_style="distributed" */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    
    wire n2319;
    wire [31:0]stack_N_397;
    
    wire stack_zc_3_1;
    wire [31:0]n1;
    
    wire Z, stack_zc_4_1, n9_c;
    wire [7:0]n1108;
    
    wire n22250, n15, stack_zc_2_1, n15_adj_460, n17, n19177, n838, 
        n2318;
    wire [4:0]n3;
    
    wire n14275, n7_c, n14, n7_adj_462, n14_adj_463;
    wire [7:0]Z_N_378;
    
    wire n14276, n14_adj_464, n15_adj_465, n19022, n16;
    wire [7:0]out_port_7__N_217;
    wire [7:0]s_N_294;
    
    wire creg_N_407, n15_adj_466, n17_adj_467, n18993, n826;
    wire [4:0]st;   // f:/home/mini-mcu/step_fpga/mcu.v(107[11:13])
    
    wire n15_adj_469, n17_adj_470, n822, n15_adj_471, n17_adj_472, 
        n818;
    wire [2:0]intr_f;   // f:/home/mini-mcu/step_fpga/mcu.v(148[11:17])
    
    wire n2312, n2317, n22288, n2316, n2315, stack_zc_1_1;
    wire [4:0]st_zc;   // f:/home/mini-mcu/step_fpga/mcu.v(119[15:20])
    
    wire n20062, n2311, jp, n22299, stack_zc_5_1, n2314, n6, n7_adj_473, 
        n16283, n8_c, n2313, n2343;
    wire [11:0]n1844;
    
    wire n2341, n2339, n2337, s_0_0, n399, s_0_1, clk_in_c_enable_16, 
        n403, s_0_2, n407, s_0_3, n411, s_0_4, n415, s_0_5, 
        n419, s_0_6, n423, s_0_7, n427, s_1_0, n431, s_1_1, 
        clk_in_c_enable_22, n435, s_1_2, n439, s_1_3, n443, s_1_4, 
        n447, s_1_5, n451, s_1_6, n455, s_1_7, n459, s_2_0, 
        n463, s_2_1, clk_in_c_enable_28, n467, s_2_2, n471, s_2_3, 
        n475, s_2_4, n479, s_2_5, n483, s_2_6, n487, s_2_7, 
        n491, s_3_0, n495, s_3_1, clk_in_c_enable_34, n499, s_3_2, 
        n503, s_3_3, n507, s_3_4, n511, s_3_5, n515, s_3_6, 
        n519, s_3_7, n523, s_4_0, n527, s_4_1, clk_in_c_enable_40, 
        n531, s_4_2, n535, s_4_3, n539, s_4_4, n543, s_4_5, 
        n547, s_4_6, n551, s_4_7, n555, s_5_0, n559, s_5_1, 
        clk_in_c_enable_46, n563, s_5_2, n567, s_5_3, n571, s_5_4, 
        n575, s_5_5, n588, s_5_6, n592, s_5_7, n596, s_6_0, 
        n600, s_6_1, clk_in_c_enable_52, n604, s_6_2, n608, s_6_3, 
        n612, s_6_4, n616, s_6_5, n620, s_6_6, n624, s_6_7, 
        n628, s_7_0, n632, s_7_1, clk_in_c_enable_58, n636, s_7_2, 
        n640, s_7_3, n645, s_7_4, n649, s_7_5, n653, s_7_6, 
        n657, s_7_7, n661, s_8_0, n665, s_8_1, clk_in_c_enable_64, 
        n669, s_8_2, n673, s_8_3, n677, s_8_4, n681, s_8_5, 
        n685, s_8_6, n689, s_8_7, n693, s_9_0, n697, s_9_1, 
        clk_in_c_enable_70, n701, s_9_2, n714, s_9_3, n718, s_9_4, 
        n722, s_9_5, n726, s_9_6, n730, s_9_7, n734, s_10_0, 
        n738, s_10_1, clk_in_c_enable_76, n742, s_10_2, n746, s_10_3, 
        n750, s_10_4, n754, s_10_5, n758, s_10_6, n762, s_10_7, 
        n766, s_11_0, n770, s_11_1, clk_in_c_enable_82, n774, s_11_2, 
        n778, s_11_3, n782, s_11_4, n786, s_11_5, n790, s_11_6, 
        n794, s_11_7, n798, s_12_0, n802, s_12_1, clk_in_c_enable_88, 
        n806, s_12_2, n810, s_12_3, n814, s_12_4, s_12_5, s_12_6, 
        s_12_7, n830, s_13_0, n834, s_13_1, clk_in_c_enable_94, 
        s_13_2, n842, s_13_3, n846, s_13_4, n850, s_13_5, n854, 
        s_13_6, n858, s_13_7, n862, s_14_0, n866, s_14_1, clk_in_c_enable_100, 
        n870, s_14_2, n874, s_14_3, n878, s_14_4, n882, s_14_5, 
        n886, s_14_6, n890, s_14_7, n894, s_15_0, n898, s_15_1, 
        clk_in_c_enable_106, n902, s_15_2, n906, s_15_3, n910, s_15_4, 
        n914, s_15_5, n918, s_15_6, n922, s_15_7, n926, n2335, 
        n15_adj_474, n17_adj_475, n19699, n19700, n7_adj_476, n15_adj_477, 
        n17_adj_478, n14261, n7_adj_479, n14_adj_480, n7_adj_481, 
        n14_adj_482;
    wire [7:0]Z_N_367;
    
    wire n14262, n15_adj_483, n17_adj_484, out_port_7__N_232, n10012;
    wire [0:0]C_N_336;
    
    wire port_id_7__N_215, n10010, n23, n23_adj_485, n23_adj_486, 
        n23_adj_487, n23_adj_488, n23_adj_489, n23_adj_490, n2333, 
        n14_adj_491, n15_adj_492, n18838, n16_adj_493, n2331, n22219, 
        n22102, n14_adj_494, n10_c, n15_adj_495, n8_adj_496, n12, 
        n18826, n13_adj_497, n15_adj_498, n17_adj_499, n18809, n2327, 
        clk_in_c_enable_109, n2730, write_strobe_N_287, n7_adj_500, 
        n14_adj_501, n14266;
    wire [17:0]n18;
    
    wire n14267, n15_adj_502, n17_adj_503, n15_adj_504, n17_adj_505, 
        n15_adj_506, n17_adj_507, n22151, n22153, n22152;
    wire [15:0]n213;
    
    wire n17550, n2325, n15_adj_508, n17_adj_509, n2329, n15_adj_510, 
        n17_adj_511, stack_zc_d0_20_0, C, n14_adj_512, n15_adj_513, 
        n18654, n16_adj_514, n22227, n22281, n13_adj_515, n13_adj_516, 
        n10_adj_517, n2322, clk_in_c_enable_115, enable_intr_flag, clk_in_c_enable_113, 
        n2320, stack_zc_d0_19_0, n22235;
    wire [7:0]port_id_7__N_200;
    
    wire n11_adj_519, n2347, n2324, n2326, n2328, n2330, n2332, 
        n2334, n2336, n2338, n2340, n2342, n2344, n2346, n22259;
    wire [7:0]n703;
    
    wire n13_adj_520, n2345, stack_zc_d0_18_0, stack_zc_d0_17_0, stack_zc_d0_16_0, 
        n15_adj_521, n17_adj_522, n18625, n15_adj_523, n17_adj_524, 
        stack_zc_d0_15_0, stack_zc_d0_14_0, stack_zc_d0_13_0, stack_zc_d0_12_0, 
        stack_zc_d0_11_0, stack_zc_d0_10_0, stack_zc_d0_9_0, stack_zc_d0_8_0, 
        stack_zc_d0_7_0, stack_zc_d0_6_0, stack_zc_d0_5_0, n15_adj_525, 
        n17_adj_526, stack_zc_d0_4_0, stack_zc_d0_3_0, stack_zc_d0_2_0, 
        stack_zc_d0_1_0, stack_zc_20_1, n22254, n12_adj_527, stack_zc_19_1, 
        stack_zc_18_1, stack_zc_17_1, stack_zc_16_1, n14_adj_528, n10_adj_529, 
        n15_adj_530, stack_zc_15_1, stack_zc_14_1, n13_adj_531;
    wire [7:0]Z_N_387;
    
    wire n22251, n14_adj_532, stack_zc_13_1, n8627, n5, n17508, 
        n20371, stack_zc_12_1, stack_zc_11_1, stack_zc_10_1, stack_zc_9_1, 
        stack_zc_8_1, n15_adj_533, n17_adj_534, stack_zc_7_1, stack_zc_6_1, 
        n15_adj_535, n17_adj_536, n22150, n22149, n22148, n15_adj_537, 
        n17_adj_538, n14_adj_539, n15_adj_540, n18321, n16_adj_541, 
        n12_adj_542, n8_adj_543, n12_adj_544, n18306, n13_adj_545, 
        n19706, n19707, n15_adj_546, n17_adj_547, n18361, n14274, 
        n15_adj_548, n17_adj_549, n15_adj_550, n17_adj_551, n15_adj_552, 
        n17_adj_553, n14286;
    wire [8:0]C_N_342;
    
    wire n15_adj_554, n17_adj_555, n15_adj_556, n17_adj_557, clk_in_c_enable_159, 
        n2755, n14_adj_558, n15_adj_559, n18286, n16_adj_560, n15_adj_561, 
        n17_adj_562, n18257;
    wire [3:0]n2634;
    
    wire n22316, n12_adj_563, n15_adj_564, n17_adj_565, n15_adj_566, 
        n17_adj_567, n15_adj_568, n17_adj_569, clk_in_c_enable_175, 
        n10021;
    wire [17:0]n1238;
    
    wire n15_adj_570, n17_adj_571, n15_adj_572, n17_adj_573, n14_adj_574, 
        n15_adj_575, n18102, n16_adj_576, n8_adj_577, n12_adj_578, 
        n18090, n13_adj_579, n12_adj_580;
    wire [17:0]pc;   // f:/home/mini-mcu/step_fpga/mcu.v(97[12:14])
    
    wire n21516, n15_adj_581, n17_adj_582, n18073, n12_adj_583, n15_adj_584, 
        n17_adj_585, n22277, n10_adj_586, n22129, n15_adj_587, n17_adj_588, 
        n15_adj_589, n17_adj_590, n15_adj_591, n17_adj_592, clk_in_c_enable_173, 
        C_N_304, clk_in_c_enable_174, Z_N_356, n23_adj_593, n15_adj_594, 
        n17_adj_595, n10_adj_596, n22228, n14_adj_597, n15_adj_598, 
        n17918, n16_adj_599, n15_adj_600, n17_adj_601, n17889, n8647, 
        n5_adj_602, n15_adj_603, n17_adj_604, n15_adj_605, n17_adj_606, 
        n15_adj_607, n17_adj_608, n19713, n19714, n7_adj_609, n22145, 
        n22147, n22146, n17366, n15_adj_610, n17_adj_611, n15_adj_612, 
        n17_adj_613, n19720, n19721, n14_adj_614, n15_adj_615, n17734, 
        n16_adj_616, n22311, n22312, n22313, n8_adj_617, n12_adj_618, 
        n17722, n13_adj_619, n12_adj_620, n15_adj_621, n17_adj_622, 
        n17705, n5_adj_623, n15_adj_624, n19727, n19728, n13_adj_625, 
        n14_adj_626, n15_adj_627, n17_adj_628, n15_adj_629, n17_adj_630, 
        n9_adj_631, n15_adj_632, n16246, n15_adj_633, n17_adj_634, 
        n15_adj_635, n17_adj_636, n19734, n19735, n15_adj_637, n17_adj_638, 
        n14_adj_639, n15_adj_640, n16_adj_641, n15_adj_642, n17_adj_643, 
        n17521, n15_adj_644, n17_adj_645, n15_adj_646, n17_adj_647, 
        n10_adj_648, n14_adj_649, n15_adj_650, n17_adj_651, n10_adj_652, 
        n14_adj_653, n11_adj_654, n13_adj_655, n14_adj_656, n13_adj_657, 
        n14_adj_658, n13_adj_659, n14_adj_660, n13_adj_661, n14_adj_662, 
        n11_adj_663, n11_adj_664, n15_adj_665, n17_adj_666, n15_adj_667, 
        n17_adj_668, n14_adj_669, n15_adj_670, n16_adj_671, n11_adj_672, 
        n11_adj_673, n17324, n20131, n12_adj_674, n17354, n13_adj_675, 
        n15_adj_676, n17_adj_677, n17337, n22144, n22143, n22142, 
        n22255, n11_adj_678, n15_adj_679, n17_adj_680, n11_adj_681, 
        n11_adj_682, n22139, n22141, n22140, n17182, n15_adj_683, 
        n17_adj_684, n11_adj_685, n11_adj_686, n11_adj_687, n22284, 
        n7746, n22307, n22236, n11_adj_688, n17140, n20199, n21794, 
        n21791, n21795, n22138, n22137, n22136, n22285, n21793, 
        n21792, n22282, n22253, n11_adj_689, n15_adj_690, n17_adj_691, 
        n11_adj_692, n160, n22117, n11_adj_693, n22133, n22135, 
        n22134, n16998, n22304, n22283, n21790, n21789, n16251, 
        n6_adj_694, n19954, n8070, n8_adj_695, n22264, n19953, n19952, 
        n19951, n13_adj_696, n22257, n14_adj_697, n10_adj_698, n22266, 
        n19950, n19949, n10_adj_699, n14_adj_700, n10_adj_701, n10_adj_702, 
        n13_adj_703, n14_adj_704, n19948, n19947, n19939, n19938, 
        n14_adj_705, n10_adj_706, n9_adj_707, n8_adj_708, n22263, 
        n14_adj_709, n10_adj_710, n19937, n14_adj_711, n10_adj_712, 
        n5_adj_713, n19936, n13_adj_714, n14_adj_715, n19935, n10_adj_716, 
        n13_adj_717, n14_adj_718, n19934, n10_adj_719, n19933, n19932, 
        n22267, n22268, n22089, n19930, n8044, n19929, n10_adj_720, 
        n19927, n19926, n21081, n6_adj_721, n7925, n8_adj_722, n15_adj_723, 
        n17_adj_724, n22094, n13_adj_725, n14_adj_726, n22099, n10_adj_727, 
        n10_adj_728, n10_adj_729;
    wire [15:0]n54;
    
    wire n10_adj_730, n13_adj_731, n5_adj_732, n10_adj_733, n14_adj_734, 
        n10_adj_735, n16349, n7946, n13_adj_736, n5_adj_737, n10_adj_738, 
        n13_adj_739, n10_adj_740, n16258, n10_adj_741, n16355, n7945, 
        n15_adj_742, n17_adj_743, n16244, n13_adj_744, n10_adj_745, 
        n7944, n22229, n11_adj_746, n16259, n16350, n10_adj_747, 
        n13_adj_748, n10_adj_749, n22246, n16727;
    wire [15:0]n151;
    
    wire n16341, n16268, n22101, n16508, n22084, n14_adj_750, n10_adj_751, 
        n15_adj_752, n55, n11_adj_753, n16532, n66, n14_adj_754, 
        n15_adj_755, n16_adj_756, n14_adj_757, n10_adj_758, n15_adj_759, 
        n14_adj_760, n10_adj_761, n15_adj_762, n11_adj_763, n56, n14413, 
        n7926, n11_adj_764, n11_adj_765, n11_adj_766, n7943, n8050, 
        n22279, n14_adj_767, n10_adj_768, n15_adj_769, n14_adj_770, 
        n10_adj_771, n15_adj_772, n14_adj_773, n10_adj_774, n15_adj_775, 
        n10_adj_776, n22093, n9_adj_777, n22085, n14_adj_778, n10_adj_779, 
        n15_adj_780, n16252, n16347, n6_adj_781, n7924, n8_adj_782, 
        n14_adj_783, n10_adj_784, n15_adj_785, n14_adj_786, n10_adj_787, 
        n15_adj_788, n14_adj_790, n10_adj_791, n15_adj_792, n14_adj_793, 
        n10_adj_794, n15_adj_795, n16269, n16338, n17_adj_796, n17153, 
        n22237, n14_adj_797, n10_adj_798, n15_adj_799, n21098, n22095, 
        n9_adj_800, n22086, n14_adj_801, n10_adj_802, n14_adj_803, 
        n10_adj_804, n14_adj_805, n10_adj_806, n16484, n22278, n14_adj_807, 
        n10_adj_808, n14_adj_809, n10_adj_810, n17_adj_811, n10_adj_812, 
        n4, n22097, n22275, n17_adj_813, n12_adj_814, n22123, n16644, 
        n22124, n22125, n16652, n20976, n9_adj_815, n17_adj_816, 
        n7923, n14_adj_817, n10_adj_818, n16956, n20317, n16331, 
        n9_adj_820, n22087, n14_adj_821, n10_adj_822, n22274, n22273, 
        n22272, n14_adj_823, n10_adj_824, n17_adj_825, n22271, n16378, 
        n14_adj_826, n10_adj_827, n22270, n22230, n11_adj_828, n22269, 
        n22132, n22131, n22130, Z_N_377, n14358, n34, n16282, 
        n17_adj_829, n16326, n6978, n8_adj_830, n14_adj_831, n10_adj_832, 
        n22222, n15_adj_833, n11_adj_834, n8789, n16253, n14_adj_835, 
        n10_adj_836;
    wire [8:0]C_N_338;
    
    wire n14422, n16245, n22231, n17906, n11804, n7052, n20, n7080, 
        n7_adj_837, n16354, n6_adj_838, n8_adj_839, n16487, n16356, 
        n19798, n19797, n19795, n14_adj_840, n15_adj_841, n16_adj_842, 
        n16389, n16_adj_843, n13_adj_844, n16391, n19794, n19792, 
        n19791, n19789, n19788, n22318, n19786, n8_adj_845, n12_adj_846, 
        n16986, n13_adj_847, n19785, n19777, n19776, n19775, n19774, 
        n19773, n22317, n16_adj_848, n16524, n14780, n19772, n19771, 
        n19770, n19768, n8_adj_849, n19767, n2, n4_adj_850, n19765, 
        n17_adj_851, n16969, n19764, n6886, n6_adj_852, n8_adj_853, 
        n19762, n19761, n17_adj_854, n19759, n19758, n19756, n19755, 
        n9164, n20152, n16685, n22082, n19753, n19752, n19750, 
        n19749, n19747, n2_adj_855, n4_adj_856, n19746, n19744, 
        n16618, n14_adj_857, n10_adj_858, n19743, n16375, n12_adj_859, 
        n12_adj_860, n5_adj_861, n14428, n17_adj_862, n10_adj_863, 
        n21531, n21796, n7628, n19, n9_adj_864, n17_adj_865, n14802, 
        n14803, n22159, n22088, n10_adj_866, n10_adj_867, n10_adj_868, 
        n10_adj_869, n17_adj_870, n20080, n10_adj_871, n11_adj_872, 
        n10_adj_873, n10_adj_874, n17_adj_875, n9_adj_876, n22165, 
        n14_adj_877, n10_adj_878, n19741, n19740, n16814, n16_adj_879, 
        n2_adj_880, n4_adj_881, n19738, n19737, n19733, n14_adj_882, 
        n10_adj_883, n19732, n6_adj_884, n8_adj_885, n19731, n14_adj_886, 
        n10_adj_887, n19730, n19726, n19725, n22232, n15_adj_888, 
        n19724, n19723, n15_adj_889, n17_adj_890, n19719, n2_adj_891, 
        n4_adj_892, n19718, n19717, n12_adj_893, n14_adj_894, n10_adj_895, 
        n12_adj_896, n19716, n14_adj_897, n10_adj_898, n14_adj_899, 
        n10_adj_900, n19712, n2_adj_901, n4_adj_902, n15_adj_903, 
        n17_adj_904, n9_adj_905, n19711, n22171, n22090, n14_adj_906, 
        n10_adj_907, n12_adj_908, n12_adj_909, n14_adj_910, n10_adj_911, 
        n14_adj_912, n10_adj_913, n6_adj_914, n8_adj_915, n19710, 
        n19709, n15_adj_916, n17_adj_917, n19705, n7066, n12_adj_918, 
        n12_adj_919, n14_adj_920, n10_adj_921, n2_adj_922, n4_adj_923, 
        n15_adj_924, n17_adj_925, n21115, n19704, n22233, n10_adj_926, 
        n2_adj_927, n4_adj_928, n14_adj_929, n10_adj_930, n19703, 
        n19702, n19698, n19697, n14_adj_931, n10_adj_932, n15_adj_933, 
        n17_adj_934, n22321, n6_adj_935, n8_adj_936, n10_adj_937, 
        n19696, n19695, n19691, n19690, n22320, n19689, n2_adj_938, 
        n4_adj_939, n19688, n13_adj_940, n19684, n19683, n2_adj_941, 
        n4_adj_942, n15_adj_943, n17_adj_944, n19682, n19681, n19673, 
        n19672, n19671, n19670, n19669, n6900, n6_adj_945, n8_adj_946, 
        n16358, n7696, n61, n16357, n19668, n2_adj_947, n4_adj_948, 
        n19667, n19666, n19658, n19657, n19656, n19655, n19654, 
        n19653, n19652, n19651, n19643, n2_adj_949, n4_adj_950, 
        n19642, n14_adj_951, n15_adj_952, n16_adj_953, n19641, n19640, 
        n13_adj_954, n13_adj_955, n1339, n1341, n21515, n9_adj_956, 
        n13_adj_957, n7094, n6_adj_958, n8_adj_959, n14_adj_960, n15_adj_961, 
        n16_adj_962, n13_adj_963, n5_adj_964, n14_adj_965, n15_adj_966, 
        n16_adj_967, n21530, n14_adj_968, n16_adj_969, n13_adj_970, 
        n2_adj_971, n4_adj_972, n14_adj_973, n15_adj_974, n16_adj_975, 
        n22177, n22091, n14_adj_976, n14_adj_977, n14_adj_978, n15_adj_979, 
        n16_adj_980, n14_adj_981, n20184, n19421, n15_adj_982, n16_adj_983, 
        n22234, n29, n24, n85, n19928, n21, n30, n19639, n14_adj_984, 
        n15_adj_985, n19390, n16_adj_986, n14_adj_987, n19206, n16_adj_988, 
        n19638, n14_adj_989, n14_adj_990, n2_adj_991, n4_adj_992, 
        n14_adj_993, n19637, n9_adj_994, n19636, n20160, n19570, 
        n6_adj_995, n8_adj_996, n22183, n22092, n14_adj_997, n10_adj_998, 
        n17339, n20077, n17362, n18075, n20164, n17213, n11_adj_999, 
        n20167, n18098, n8773, n14_adj_1000, n10_adj_1001, n21132, 
        n14_adj_1002, n10_adj_1003, n14_adj_1004, n10_adj_1005, n19628, 
        n19627, n14_adj_1006, n10_adj_1007, n14_adj_1008, n10_adj_1009, 
        n9_adj_1010, n2_adj_1011, n4_adj_1012, n18811, n22189, n14_adj_1013, 
        n11_adj_1014, n19626, n19625, n2_adj_1015, n4_adj_1016, n11_adj_1017, 
        n19624, n19623, n14_adj_1018, n19622, n19621, n2_adj_1019, 
        n4_adj_1020, n19613, n14_adj_1021, n19612, n19611, n19610, 
        n22324, n14_adj_1022, n19609, n19608, n11_adj_1023, n14_adj_1024, 
        n15_adj_1025, n16_adj_1026, n19607, n19606, n14_adj_1027, 
        n19598, n19597, n19596, n11_adj_1028, n19595, n19594, n11_adj_1029, 
        n19593, n19592, n19591, n19583, n20203, n17949, n19582, 
        n19581, n19580, n14_adj_1030, n19579, n19578, n19577, n19576, 
        n9_adj_1031, n22195, n22096, n14_adj_1032, n10_adj_1033, n14_adj_1034, 
        n10_adj_1035, n11_adj_1036, n20914, n14_adj_1037, n10_adj_1038, 
        n21529, n22323, n21187, n4_adj_1039, n4_adj_1040, n63_adj_1041, 
        n10_adj_1042, n14285, n14_adj_1043, n10_adj_1044, n14_adj_1045, 
        n10_adj_1046, n14_adj_1047, n10_adj_1048, n14284, n11_adj_1049, 
        n9_adj_1050, n14283, n20324, n18834, n22213, n22098, n14_adj_1051, 
        n12_adj_1052, n14_adj_1053, n20358, n18685, n19547, n14_adj_1054, 
        n22119, n14_adj_1055, n14_adj_1056, n22327, n14_adj_1057, 
        n22122, n14_adj_1058, n10_adj_1059, n15_adj_1060, n14_adj_1061, 
        n10_adj_1062, n15_adj_1063, n22238, n12_adj_1064, n12_adj_1065, 
        n12_adj_1066, n22100, n14_adj_1067, n10_adj_1068, n15_adj_1069, 
        n22309, n12_adj_1070, n22326, n10_adj_1073, n12_adj_1074, 
        n12_adj_1075, n14_adj_1076, n10_adj_1077, n15_adj_1078, n14_adj_1079, 
        n10_adj_1080, n15_adj_1081, n14_adj_1082, n15_adj_1083, n16_adj_1084, 
        n14_adj_1085, n10_adj_1086, n15_adj_1087, n22116, n14_adj_1088, 
        n10_adj_1089, n15_adj_1090, n5_adj_1091, n15_adj_1092, n14_adj_1093, 
        n10_adj_1094, n15_adj_1095, n10_adj_1096, n10_adj_1097, n14_adj_1098, 
        n15_adj_1099, n22239, n10_adj_1100, n14_adj_1101, n15_adj_1102, 
        n16_adj_1103, n17_adj_1104, n14_adj_1105, n15_adj_1106, n20955, 
        n10_adj_1107, n16_adj_1108, n17_adj_1109, n14_adj_1110, n15_adj_1111, 
        n16_adj_1112, n17_adj_1113, n16_adj_1114, n17_adj_1115, n9_adj_1116, 
        n16_adj_1117, n17_adj_1118, n21170, n14263, n16_adj_1119, 
        n17_adj_1120, n17370, n18106, n13_adj_1121, n18842, n21186, 
        n13_adj_1124, n13_adj_1125, n22214, n22218, n19164, n20268, 
        n13_adj_1128, n20349, n13_adj_1129, n22217, n22216, n22215, 
        n13_adj_1130, n20366, n14_adj_1131, n16_adj_1132, n17002, 
        n17738, n18474, n22240, n20089, n14265, n22083, n19210, 
        n10_adj_1133, n22308, n22245, n11_adj_1136, n20144, n11_adj_1137, 
        n22118, n11_adj_1138, n11_adj_1139, n11_adj_1140, n22261, 
        n22205, n17186, n11_adj_1141, n19394, n15_adj_1142, n16_adj_1143, 
        n11_adj_1144, n11_adj_1145, n20177, n17922, n18658, n22248, 
        n18274, n12_adj_1146, n12_adj_1147, n5_adj_1148, n12_adj_1149, 
        n16818, n1124, n20258, n16122, n103, n16123, n12_adj_1150, 
        n12_adj_1151, n20312, n12_adj_1152, n17554, n12_adj_1153, 
        n12_adj_1154, n18290, n19026;
    wire [17:0]n1194;
    
    wire n5_adj_1155, n2323;
    wire [11:0]n1742;
    
    wire n14264, n20074, n14459, n22252, n10_adj_1156, n10_adj_1157, 
        n12_adj_1158, n5_adj_1159, n13_adj_1160, n14_adj_1161, n15_adj_1162, 
        n16_adj_1163, n12_adj_1164, n12_adj_1165, n13_adj_1166, n13_adj_1167, 
        n12_adj_1168, n12_adj_1169, n13_adj_1170, n12_adj_1171, n13_adj_1172, 
        n13_adj_1173, n5_adj_1174, n9_adj_1175, n15_adj_1176, n14414, 
        n10_adj_1177, n13_adj_1178, n11_adj_1179, n14_adj_1180, n15_adj_1181, 
        n16_adj_1182, n5_adj_1183, n13_adj_1184, n13_adj_1185, n11_adj_1186, 
        n13_adj_1187, n11_adj_1188, n11_adj_1189, n13_adj_1190, n11_adj_1191, 
        n11_adj_1192, n13_adj_1193, n11_adj_1194, n11_adj_1195, n22258, 
        n12_adj_1196, n20194, n19361, n14270, n20305, n10_adj_1197, 
        n21201, n20384, n17397, n20128, n18282, n5_adj_1198, n1384;
    wire [0:0]C_N_351;
    
    wire n77, n17523, n20354, n17546, n20155, n18133, n20292, 
        n19018, n18259, n19793, n14_adj_1199, n20321, n18869, n12_adj_1200, 
        n18995, n12_adj_1201, n19787, n12_adj_1202, n12_adj_1203, 
        n12_adj_1204, n12_adj_1205, n5_adj_1206, n10_adj_1207, n10_adj_1208, 
        n13_adj_1209, n13_adj_1210, n13_adj_1211, n13_adj_1212, n13_adj_1213, 
        n13_adj_1214, n14_adj_1215, n15_adj_1216, n19574, n16_adj_1217, 
        n19633, n19634, n20302, n16994, n17707, n20375, n16845, 
        n20297, n17730, n18363, n20346, n17581, n14281, n20382, 
        n18466, n19179, n20095, n18317, n20263, n19202, n16971, 
        n11_adj_1218, n20285, n19053, n21226, n11_adj_1219, n11_adj_1220, 
        n11_adj_1221, n11_adj_1222, n11_adj_1223, n11_adj_1224, n11_adj_1225, 
        n16522, n11_adj_1226, n11_adj_1227, n18642, n16_adj_1228, 
        n16_adj_1229, n17_adj_1230, n12_adj_1231, n22249, n12_adj_1232, 
        n16_adj_1233, n17_adj_1234, n16_adj_1235, n17_adj_1236, n16_adj_1237, 
        n17_adj_1238, n6928, n16792, n12_adj_1240, n16_adj_1241, n17_adj_1242, 
        n12_adj_1243, n12_adj_1244, n12_adj_1245, n12_adj_1246, n12_adj_1247, 
        n19754, n5_adj_1248, n10_adj_1249, n10_adj_1250, n13_adj_1251, 
        n13_adj_1252, n19796, n13_adj_1253, n13_adj_1254, n13_adj_1255, 
        n13_adj_1256, n22114, n22115, n19532, n20170, n22108, n22112, 
        n22113, n10_adj_1257, n6914, n11916, n22221, n14280, n22276, 
        n11_adj_1258, n11_adj_1259, n22120, n22121, n19348, n11_adj_1260, 
        n14279, n22107, n22110, n22111, n11_adj_1261, n10_adj_1262, 
        n11_adj_1263, n16558, n22291, n11_adj_1264, n16409, n21644, 
        n11_adj_1265, n11_adj_1266, n22300, n12_adj_1267, n10_adj_1268, 
        n10_adj_1269, n21255, n22211, n22212, n22163, n22187, n22126, 
        n16672, n22128, n22127, n16_adj_1270, n22169, n22193, n16_adj_1271, 
        n22175, n14278, n16_adj_1272, n22305, n16_adj_1273, n16_adj_1274, 
        n16_adj_1275, n22157, n22181, n11_adj_1276, n22306, n12_adj_1277, 
        n11_adj_1278, n19742, n12_adj_1279, n12_adj_1280, n12_adj_1281, 
        n19748, n11_adj_1282, n48, n12_adj_1283, n12_adj_1284, n11_adj_1285, 
        n11_adj_1286, n10_adj_1287, n10_adj_1288, n8_adj_1289, n13_adj_1290, 
        n13_adj_1291, n13_adj_1292, n13_adj_1293, n13_adj_1294, n13_adj_1295, 
        n11_adj_1296, n22103, n22247, n16_adj_1297, n17_adj_1298, 
        n16_adj_1299, n17_adj_1300, n16_adj_1301, n17_adj_1302, n22104, 
        n22105, n11_adj_1303, n11_adj_1304, n19545, n16_adj_1305, 
        n17_adj_1306, n16_adj_1307, n17_adj_1308, n22197, n16_adj_1309, 
        n17_adj_1310, n22199, n22200, n22201, n22242, n16_adj_1311, 
        n22202, n16_adj_1312, n16_adj_1313, n16_adj_1314, n16_adj_1315, 
        n16_adj_1316, n22280, n22203, n22204, n12_adj_1317, n16_adj_1318, 
        n16_adj_1319, n16_adj_1320, n16_adj_1321, n22206, n16_adj_1322, 
        n16662, n16800, n22196, n16_adj_1323, n16_adj_1324, n16_adj_1325, 
        n16_adj_1326, n16_adj_1327, n16_adj_1328, n16_adj_1329, n22209, 
        n12_adj_1330, n18980, n22210, n22208, n22207, n16_adj_1331, 
        n16_adj_1332, n16_adj_1333, n16_adj_1334, n16_adj_1335, n16_adj_1336, 
        n12_adj_1337, n22244, n16_adj_1338, n16_adj_1339, n16_adj_1340, 
        n16_adj_1341, n12_adj_1342, n12_adj_1343, n16_adj_1344, n16_adj_1345, 
        n19961, n12_adj_1346, n16701, n10_adj_1347, n16_adj_1348, 
        n10_adj_1349, n10_adj_1350, n10_adj_1351, n16_adj_1352, n12_adj_1353, 
        n16_adj_1354, n16_adj_1355, n16_adj_1356, n16_adj_1357, n16_adj_1358, 
        n16_adj_1359, n17_adj_1360;
    wire [15:0]n346;
    
    wire n17_adj_1361, n16_adj_1362, n14269, n16_adj_1363, n16_adj_1364, 
        n16_adj_1365, n17_adj_1366, n17_adj_1367, n17_adj_1368, n17_adj_1369, 
        n16590, n22243, n17_adj_1370, n10_adj_1371, n17_adj_1372, 
        n17_adj_1373, n17_adj_1374, n22260, n16_adj_1375, n22325, 
        n16574, n17_adj_1376, n10_adj_1377, n17_adj_1378, n17_adj_1379, 
        n13_adj_1380, n17_adj_1381, n22198, n17_adj_1382, n16_adj_1383, 
        n13_adj_1384, n17_adj_1385, n17_adj_1386, n13_adj_1387, n17_adj_1388, 
        n17_adj_1389, n13_adj_1390, n17_adj_1391, n22256, n16_adj_1392, 
        n17_adj_1393, n13_adj_1394, n17_adj_1395, n13_adj_1396, n17_adj_1397, 
        n17_adj_1398, n22241, n17_adj_1399, n16364, n16_adj_1400, 
        n16_adj_1401, n19766, n16_adj_1402, n19760, n19663, n19664, 
        n19618, n19619, n16_adj_1403, n19588, n19589, n19603, n19604, 
        n19648, n19649, n19782, n19783, n11_adj_1404, n11_adj_1405, 
        n11_adj_1406, n22194, n11_adj_1407, n6_adj_1408, n11_adj_1409, 
        n11_adj_1410, n11_adj_1411, n11_adj_1412, n11_adj_1413, n11_adj_1414, 
        n11_adj_1415, n18796, n22192, n22191, n22190, n8_adj_1416, 
        n14_adj_1417, n16636, n11_adj_1418, n50, n16_adj_1419, n11_adj_1420, 
        n22188, n16810, n16_adj_1421, n16_adj_1422;
    wire [3:0]n2641;
    
    wire n16_adj_1423, n11_adj_1424, n16_adj_1425, n16_adj_1426, n19010, 
        n12_adj_1427, n12_adj_1428, n18612, n22186, n22185, n22184, 
        n5_adj_1429, n4_adj_1430, n11_adj_1431, n11_adj_1432, n12_adj_1433, 
        n12_adj_1434, n12_adj_1435, n11_adj_1436, n12_adj_1437, n12_adj_1438, 
        n17170, n11_adj_1439, n12_adj_1440, n12_adj_1441, n12_adj_1442, 
        n11_adj_1443, n19363, n12_adj_1444, n22182, n11_adj_1445, 
        n6_adj_1446, n12_adj_1447, n18368, n22180, n22179, n22178, 
        n10_adj_1448, n22176, n12_adj_1449, n10_adj_1450, n18244, 
        n22174, n22173, n22172, n13_adj_1451, n13_adj_1452, n22287, 
        n8_adj_1453, n17_adj_1454, n15_adj_1455, n11_adj_1456, n9_adj_1457, 
        n22322, n7_adj_1458, n21532, n13_adj_1459, n13_adj_1460, n12_adj_1461, 
        n18627, n13_adj_1462, n12_adj_1463, n22170, n6_adj_1464, n12_adj_1465, 
        n9_adj_1466, n12_adj_1467, n12_adj_1468, n22319, n105, n22328, 
        n13_adj_1469, n10_adj_1470, n18060, n22106, n22168, n22167, 
        n22166, n75, n71, n14425, n53, n16239;
    wire [0:0]C_N_352;
    
    wire n19946, n22, n19931, n22298, n10_adj_1471, n17891, n11_adj_1472, 
        n13_adj_1473, n13_adj_1474, n16802, n6_adj_1475, n11196, n11_adj_1476, 
        n12_adj_1477, n11_adj_1478, n11_adj_1479, n11_adj_1480, n12_adj_1481, 
        n11_adj_1482, n11_adj_1483, n11_adj_1484, n12_adj_1485, n13_adj_1486, 
        n13_adj_1487, n13_adj_1488, n11_adj_1489, n12_adj_1490, n14423, 
        n83_adj_1491, n64_adj_1492, n12_adj_1493, n16_adj_1494, n16236, 
        n14417, n16596, n12_adj_1495, n16_adj_1496, n11_adj_1497, 
        n17155, n16_adj_1498, n16_adj_1499, n16_adj_1500, n16_adj_1501, 
        n19678, n19679, n13_adj_1502, n12_adj_1503, n14_adj_1504, 
        n15_adj_1505, n14_adj_1506, n22164, n12_adj_1507, n12_adj_1508, 
        n17876, n22162, n22161, n22160, n12_adj_1509, n14_adj_1510, 
        n15_adj_1511, n22158, n6_adj_1512, n17_adj_1513, n12182, n12_adj_1514, 
        n12_adj_1515, n12_adj_1516, n12_adj_1517, n22156, n22155, 
        n22154, n17692, n12_adj_1518, n12_adj_1519, n14_adj_1520, 
        n15_adj_1521, n19194, n12_adj_1522, n12_adj_1523, n12_adj_1524, 
        n10_adj_1525, n22225, n22224, n22226, n16622, n20344, n14_adj_1526, 
        n22220, n16_adj_1527, n12_adj_1528, n13_adj_1529, n13_adj_1530, 
        n13_adj_1531, n13_adj_1532, n16_adj_1533, n13_adj_1534, n16_adj_1535, 
        n16518, n4_adj_1536, n16520, n11_adj_1537, n12_adj_1538, n16_adj_1539, 
        n13_adj_1540, n10_adj_1541, n19556, n11_adj_1542, n12_adj_1543, 
        n16_adj_1544, n10_adj_1545, n16_adj_1546, n16_adj_1547, n19403, 
        n21001, n10_adj_1548, n14_adj_1549, n16_adj_1550, n19372, 
        n20189, n16_adj_1551, n16_adj_1552, n13_adj_1553, n16_adj_1554, 
        n13_adj_1555, n16_adj_1556, n11_adj_1557, n12_adj_1558, n19219, 
        n20251, n11_adj_1559, n12_adj_1560, n13_adj_1561, n14268, 
        n13_adj_1562, n11_adj_1563, n19188, n13_adj_1564, n11_adj_1565, 
        n13_adj_1566, n19035, n11_adj_1567, n11_adj_1568;
    wire [7:0]n2055;
    
    wire n22315, n22314, n21018, n11_adj_1569, n12_adj_1570, n11_adj_1571, 
        n12_adj_1572, n19004, n11_adj_1573, n18851, n11_adj_1574, 
        n21062, n11_adj_1575, n11_adj_1576, n18820, n11_adj_1577, 
        n12_adj_1578, n18667, n22223, n11_adj_1579, n12_adj_1580, 
        n10_adj_1581, n12_adj_1582, n18636, n20361, n18483, n20377, 
        n14277, n16633, n18452, n11_adj_1583, n6_adj_1584, n18299, 
        n11_adj_1585, n18268, n19378, n17538, n18115, n12_adj_1586, 
        n11_adj_1587, n12_adj_1588, n12_adj_1589, n18084, n11_adj_1590, 
        n12_adj_1591, n17_adj_1592, n17931, n17_adj_1593, n11_adj_1594, 
        n12_adj_1595, n12_adj_1596, n11_adj_1597, n12_adj_1598, n17900, 
        n20231, n12_adj_1599, n21035, n12_adj_1600, n12_adj_1601, 
        n17747, n20287, n4_adj_1602, n19562, n17716, n17563, n10_adj_1603, 
        n10_adj_1604, n13_adj_1605, n17532, n13_adj_1606, n13_adj_1607, 
        n17379, n13_adj_1608, n13_adj_1609, n13_adj_1610, n17_adj_1611, 
        n5_adj_1612, n17_adj_1613, n15_adj_1614, n17348, n13_adj_1615, 
        n17195, n13_adj_1616, n10_adj_1617, n13_adj_1618, n17164, 
        n20182, n13_adj_1619, n16_adj_1620, n13_adj_1621, n13_adj_1622, 
        n19237, n13_adj_1623, n16_adj_1624, n19386, n13_adj_1625, 
        n13_adj_1626, n13_adj_1627, n16_adj_1628, n13_adj_1629, n13_adj_1630, 
        n11_adj_1631, n19584, n19585, n19586, n19587, n19599, n19600, 
        n13_adj_1632, n19601, n19602, n19614, n19615, n13_adj_1633, 
        n13_adj_1634, n18650, n19616, n19617, n19629, n19630, n19631, 
        n19632, n13_adj_1635, n18501, n19644, n19645, n19646, n19647, 
        n19659, n19660, n11_adj_1636, n19661, n19662, n13_adj_1637, 
        n19674, n19675, n19676, n19677, n13_adj_1638, n19778, n19779, 
        n13_adj_1639, n19780, n19781, n13_adj_1640, n13_adj_1641, 
        n17914, n13_adj_1642, n17765, n13_adj_1643, n13_adj_1644, 
        n13_adj_1645, n12_adj_1646, n13_adj_1647, n17_adj_1648, n13_adj_1649, 
        n13_adj_1650, n17178, n17_adj_1651, n13_adj_1652, n17029, 
        n13_adj_1653, n13_adj_1654, n13_adj_1655, n58, n10_adj_1656, 
        n20289, n17011, n19685, n19686, n19692, n19693, n16980, 
        n14_adj_1657, n16827, n19944, n19945, n19959, n19960, n19940, 
        n19941, n19942, n19943, n19955, n19956, n19957, n19958;
    
    FD1S3AX stack_1008 (.D(stack_N_397[4]), .CK(clk_in_c), .Q(n2319));   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam stack_1008.GSR = "ENABLED";
    FD1P3AX i24_25 (.D(Z), .SP(n1[3]), .CK(clk_in_c), .Q(stack_zc_3_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i24_25.GSR = "ENABLED";
    FD1P3AX i30_31 (.D(Z), .SP(n1[4]), .CK(clk_in_c), .Q(stack_zc_4_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i30_31.GSR = "ENABLED";
    LUT4 PrioSelect_105_i15_3_lut_4_lut_4_lut (.A(n11714), .B(n9_c), .C(n1108[7]), 
         .D(n22250), .Z(n15)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_105_i15_3_lut_4_lut_4_lut.init = 16'hccd8;
    FD1P3AX i18_19 (.D(Z), .SP(n1[2]), .CK(clk_in_c), .Q(stack_zc_2_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i18_19.GSR = "ENABLED";
    PFUMX PrioSelect_497_i19 (.BLUT(n15_adj_460), .ALUT(n17), .C0(n19177), 
          .Z(n838)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1S3AX stack_1007 (.D(n3[3]), .CK(clk_in_c), .Q(n2318));   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam stack_1007.GSR = "ENABLED";
    CCU2D add_412_5 (.A0(instruction[3]), .B0(instruction[11]), .C0(n7_c), 
          .D0(n14), .A1(instruction[4]), .B1(instruction[11]), .C1(n7_adj_462), 
          .D1(n14_adj_463), .CIN(n14275), .COUT(n14276), .S0(Z_N_378[3]), 
          .S1(Z_N_378[4]));   // f:/home/mini-mcu/step_fpga/mcu.v(275[74:85])
    defparam add_412_5.INIT0 = 16'ha965;
    defparam add_412_5.INIT1 = 16'ha965;
    defparam add_412_5.INJECT1_0 = "NO";
    defparam add_412_5.INJECT1_1 = "NO";
    PFUMX PrioSelect_489_i16 (.BLUT(n14_adj_464), .ALUT(n15_adj_465), .C0(n19022), 
          .Z(n16)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    SPR16X4C creg1 (.DI0(out_port_7__N_217[0]), .DI1(s_N_294[1]), .DI2(s_N_294[2]), 
            .DI3(s_N_294[3]), .AD0(instruction[0]), .AD1(instruction[1]), 
            .AD2(instruction[2]), .AD3(instruction[3]), .CK(clk_in_c), 
            .WRE(creg_N_407), .DO0(n1108[0]), .DO1(n1108[1]), .DO2(n1108[2]), 
            .DO3(n1108[3]));
    defparam creg1.initval = "0x0000000000000000";
    PFUMX PrioSelect_485_i19 (.BLUT(n15_adj_466), .ALUT(n17_adj_467), .C0(n18993), 
          .Z(n826)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1S3AX st__i0 (.D(n3[0]), .CK(clk_in_c), .Q(st[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam st__i0.GSR = "ENABLED";
    PFUMX PrioSelect_481_i19 (.BLUT(n15_adj_469), .ALUT(n17_adj_470), .C0(n18993), 
          .Z(n822)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_477_i19 (.BLUT(n15_adj_471), .ALUT(n17_adj_472), .C0(n18993), 
          .Z(n818)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1S3IX intr_f__i0 (.D(interrupt), .CK(clk_in_c), .CD(n22301), .Q(intr_f[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(154[8] 157[4])
    defparam intr_f__i0.GSR = "ENABLED";
    FD1S3AX stack_1001 (.D(n3[0]), .CK(clk_in_c), .Q(n2312));   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam stack_1001.GSR = "ENABLED";
    FD1S3AX stack_1006 (.D(n22288), .CK(clk_in_c), .Q(n2317));   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam stack_1006.GSR = "ENABLED";
    FD1S3AX stack_1005 (.D(n3[2]), .CK(clk_in_c), .Q(n2316));   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam stack_1005.GSR = "ENABLED";
    FD1S3AX stack_1004 (.D(stack_N_397[2]), .CK(clk_in_c), .Q(n2315));   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam stack_1004.GSR = "ENABLED";
    FD1P3AX i12_13 (.D(Z), .SP(n1[1]), .CK(clk_in_c), .Q(stack_zc_1_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i12_13.GSR = "ENABLED";
    FD1S3IX st_zc__i0 (.D(n20062), .CK(clk_in_c), .CD(n22301), .Q(st_zc[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam st_zc__i0.GSR = "ENABLED";
    FD1S3AX stack_1000 (.D(stack_N_397[0]), .CK(clk_in_c), .Q(n2311));   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam stack_1000.GSR = "ENABLED";
    FD1S3JX jp_503 (.D(n22299), .CK(clk_in_c), .PD(n22301), .Q(jp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam jp_503.GSR = "ENABLED";
    FD1P3AX i36_37 (.D(Z), .SP(n1[5]), .CK(clk_in_c), .Q(stack_zc_5_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i36_37.GSR = "ENABLED";
    FD1S3AX stack_1003 (.D(n3[1]), .CK(clk_in_c), .Q(n2314));   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam stack_1003.GSR = "ENABLED";
    LUT4 PrioSelect_201_i8_4_lut (.A(n6), .B(n7_adj_473), .C(n16283), 
         .D(n16290), .Z(n8_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_201_i8_4_lut.init = 16'hcfca;
    FD1S3AX stack_1002 (.D(stack_N_397[1]), .CK(clk_in_c), .Q(n2313));   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam stack_1002.GSR = "ENABLED";
    FD1S3AX stack_1022 (.D(n1844[9]), .CK(clk_in_c), .Q(n2343));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1022.GSR = "ENABLED";
    FD1S3AX stack_1021 (.D(n1844[8]), .CK(clk_in_c), .Q(n2341));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1021.GSR = "ENABLED";
    FD1S3AX stack_1020 (.D(n1844[7]), .CK(clk_in_c), .Q(n2339));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1020.GSR = "ENABLED";
    FD1S3AX stack_1019 (.D(n1844[6]), .CK(clk_in_c), .Q(n2337));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1019.GSR = "ENABLED";
    FD1S3AX s_0_0_c (.D(n399), .CK(clk_in_c), .Q(s_0_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_0_0_c.GSR = "ENABLED";
    FD1P3AX s_0_1_c (.D(n403), .SP(clk_in_c_enable_16), .CK(clk_in_c), 
            .Q(s_0_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_0_1_c.GSR = "ENABLED";
    FD1P3AX s_0_2_c (.D(n407), .SP(clk_in_c_enable_16), .CK(clk_in_c), 
            .Q(s_0_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_0_2_c.GSR = "ENABLED";
    FD1P3AX s_0_3_c (.D(n411), .SP(clk_in_c_enable_16), .CK(clk_in_c), 
            .Q(s_0_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_0_3_c.GSR = "ENABLED";
    FD1P3AX s_0_4_c (.D(n415), .SP(clk_in_c_enable_16), .CK(clk_in_c), 
            .Q(s_0_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_0_4_c.GSR = "ENABLED";
    FD1P3AX s_0_5_c (.D(n419), .SP(clk_in_c_enable_16), .CK(clk_in_c), 
            .Q(s_0_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_0_5_c.GSR = "ENABLED";
    FD1P3AX s_0_6_c (.D(n423), .SP(clk_in_c_enable_16), .CK(clk_in_c), 
            .Q(s_0_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_0_6_c.GSR = "ENABLED";
    FD1S3AX s_0_7_c (.D(n427), .CK(clk_in_c), .Q(s_0_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_0_7_c.GSR = "ENABLED";
    FD1S3AX s_1_0_c (.D(n431), .CK(clk_in_c), .Q(s_1_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_1_0_c.GSR = "ENABLED";
    FD1P3AX s_1_1_c (.D(n435), .SP(clk_in_c_enable_22), .CK(clk_in_c), 
            .Q(s_1_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_1_1_c.GSR = "ENABLED";
    FD1P3AX s_1_2_c (.D(n439), .SP(clk_in_c_enable_22), .CK(clk_in_c), 
            .Q(s_1_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_1_2_c.GSR = "ENABLED";
    FD1P3AX s_1_3_c (.D(n443), .SP(clk_in_c_enable_22), .CK(clk_in_c), 
            .Q(s_1_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_1_3_c.GSR = "ENABLED";
    FD1P3AX s_1_4_c (.D(n447), .SP(clk_in_c_enable_22), .CK(clk_in_c), 
            .Q(s_1_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_1_4_c.GSR = "ENABLED";
    FD1P3AX s_1_5_c (.D(n451), .SP(clk_in_c_enable_22), .CK(clk_in_c), 
            .Q(s_1_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_1_5_c.GSR = "ENABLED";
    FD1P3AX s_1_6_c (.D(n455), .SP(clk_in_c_enable_22), .CK(clk_in_c), 
            .Q(s_1_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_1_6_c.GSR = "ENABLED";
    FD1S3AX s_1_7_c (.D(n459), .CK(clk_in_c), .Q(s_1_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_1_7_c.GSR = "ENABLED";
    FD1S3AX s_2_0_c (.D(n463), .CK(clk_in_c), .Q(s_2_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_2_0_c.GSR = "ENABLED";
    FD1P3AX s_2_1_c (.D(n467), .SP(clk_in_c_enable_28), .CK(clk_in_c), 
            .Q(s_2_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_2_1_c.GSR = "ENABLED";
    FD1P3AX s_2_2_c (.D(n471), .SP(clk_in_c_enable_28), .CK(clk_in_c), 
            .Q(s_2_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_2_2_c.GSR = "ENABLED";
    FD1P3AX s_2_3_c (.D(n475), .SP(clk_in_c_enable_28), .CK(clk_in_c), 
            .Q(s_2_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_2_3_c.GSR = "ENABLED";
    FD1P3AX s_2_4_c (.D(n479), .SP(clk_in_c_enable_28), .CK(clk_in_c), 
            .Q(s_2_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_2_4_c.GSR = "ENABLED";
    FD1P3AX s_2_5_c (.D(n483), .SP(clk_in_c_enable_28), .CK(clk_in_c), 
            .Q(s_2_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_2_5_c.GSR = "ENABLED";
    FD1P3AX s_2_6_c (.D(n487), .SP(clk_in_c_enable_28), .CK(clk_in_c), 
            .Q(s_2_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_2_6_c.GSR = "ENABLED";
    FD1S3AX s_2_7_c (.D(n491), .CK(clk_in_c), .Q(s_2_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_2_7_c.GSR = "ENABLED";
    FD1S3AX s_3_0_c (.D(n495), .CK(clk_in_c), .Q(s_3_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_3_0_c.GSR = "ENABLED";
    FD1P3AX s_3_1_c (.D(n499), .SP(clk_in_c_enable_34), .CK(clk_in_c), 
            .Q(s_3_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_3_1_c.GSR = "ENABLED";
    FD1P3AX s_3_2_c (.D(n503), .SP(clk_in_c_enable_34), .CK(clk_in_c), 
            .Q(s_3_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_3_2_c.GSR = "ENABLED";
    FD1P3AX s_3_3_c (.D(n507), .SP(clk_in_c_enable_34), .CK(clk_in_c), 
            .Q(s_3_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_3_3_c.GSR = "ENABLED";
    FD1P3AX s_3_4_c (.D(n511), .SP(clk_in_c_enable_34), .CK(clk_in_c), 
            .Q(s_3_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_3_4_c.GSR = "ENABLED";
    FD1P3AX s_3_5_c (.D(n515), .SP(clk_in_c_enable_34), .CK(clk_in_c), 
            .Q(s_3_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_3_5_c.GSR = "ENABLED";
    FD1P3AX s_3_6_c (.D(n519), .SP(clk_in_c_enable_34), .CK(clk_in_c), 
            .Q(s_3_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_3_6_c.GSR = "ENABLED";
    FD1S3AX s_3_7_c (.D(n523), .CK(clk_in_c), .Q(s_3_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_3_7_c.GSR = "ENABLED";
    FD1S3AX s_4_0_c (.D(n527), .CK(clk_in_c), .Q(s_4_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_4_0_c.GSR = "ENABLED";
    FD1P3AX s_4_1_c (.D(n531), .SP(clk_in_c_enable_40), .CK(clk_in_c), 
            .Q(s_4_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_4_1_c.GSR = "ENABLED";
    FD1P3AX s_4_2_c (.D(n535), .SP(clk_in_c_enable_40), .CK(clk_in_c), 
            .Q(s_4_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_4_2_c.GSR = "ENABLED";
    FD1P3AX s_4_3_c (.D(n539), .SP(clk_in_c_enable_40), .CK(clk_in_c), 
            .Q(s_4_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_4_3_c.GSR = "ENABLED";
    FD1P3AX s_4_4_c (.D(n543), .SP(clk_in_c_enable_40), .CK(clk_in_c), 
            .Q(s_4_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_4_4_c.GSR = "ENABLED";
    FD1P3AX s_4_5_c (.D(n547), .SP(clk_in_c_enable_40), .CK(clk_in_c), 
            .Q(s_4_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_4_5_c.GSR = "ENABLED";
    FD1P3AX s_4_6_c (.D(n551), .SP(clk_in_c_enable_40), .CK(clk_in_c), 
            .Q(s_4_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_4_6_c.GSR = "ENABLED";
    FD1S3AX s_4_7_c (.D(n555), .CK(clk_in_c), .Q(s_4_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_4_7_c.GSR = "ENABLED";
    FD1S3AX s_5_0_c (.D(n559), .CK(clk_in_c), .Q(s_5_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_5_0_c.GSR = "ENABLED";
    FD1P3AX s_5_1_c (.D(n563), .SP(clk_in_c_enable_46), .CK(clk_in_c), 
            .Q(s_5_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_5_1_c.GSR = "ENABLED";
    FD1P3AX s_5_2_c (.D(n567), .SP(clk_in_c_enable_46), .CK(clk_in_c), 
            .Q(s_5_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_5_2_c.GSR = "ENABLED";
    FD1P3AX s_5_3_c (.D(n571), .SP(clk_in_c_enable_46), .CK(clk_in_c), 
            .Q(s_5_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_5_3_c.GSR = "ENABLED";
    FD1P3AX s_5_4_c (.D(n575), .SP(clk_in_c_enable_46), .CK(clk_in_c), 
            .Q(s_5_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_5_4_c.GSR = "ENABLED";
    FD1P3AX s_5_5_c (.D(n588), .SP(clk_in_c_enable_46), .CK(clk_in_c), 
            .Q(s_5_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_5_5_c.GSR = "ENABLED";
    FD1P3AX s_5_6_c (.D(n592), .SP(clk_in_c_enable_46), .CK(clk_in_c), 
            .Q(s_5_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_5_6_c.GSR = "ENABLED";
    FD1S3AX s_5_7_c (.D(n596), .CK(clk_in_c), .Q(s_5_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_5_7_c.GSR = "ENABLED";
    FD1S3AX s_6_0_c (.D(n600), .CK(clk_in_c), .Q(s_6_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_6_0_c.GSR = "ENABLED";
    FD1P3AX s_6_1_c (.D(n604), .SP(clk_in_c_enable_52), .CK(clk_in_c), 
            .Q(s_6_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_6_1_c.GSR = "ENABLED";
    FD1P3AX s_6_2_c (.D(n608), .SP(clk_in_c_enable_52), .CK(clk_in_c), 
            .Q(s_6_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_6_2_c.GSR = "ENABLED";
    FD1P3AX s_6_3_c (.D(n612), .SP(clk_in_c_enable_52), .CK(clk_in_c), 
            .Q(s_6_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_6_3_c.GSR = "ENABLED";
    FD1P3AX s_6_4_c (.D(n616), .SP(clk_in_c_enable_52), .CK(clk_in_c), 
            .Q(s_6_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_6_4_c.GSR = "ENABLED";
    FD1P3AX s_6_5_c (.D(n620), .SP(clk_in_c_enable_52), .CK(clk_in_c), 
            .Q(s_6_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_6_5_c.GSR = "ENABLED";
    FD1P3AX s_6_6_c (.D(n624), .SP(clk_in_c_enable_52), .CK(clk_in_c), 
            .Q(s_6_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_6_6_c.GSR = "ENABLED";
    FD1S3AX s_6_7_c (.D(n628), .CK(clk_in_c), .Q(s_6_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_6_7_c.GSR = "ENABLED";
    FD1S3AX s_7_0_c (.D(n632), .CK(clk_in_c), .Q(s_7_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_7_0_c.GSR = "ENABLED";
    FD1P3AX s_7_1_c (.D(n636), .SP(clk_in_c_enable_58), .CK(clk_in_c), 
            .Q(s_7_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_7_1_c.GSR = "ENABLED";
    FD1P3AX s_7_2_c (.D(n640), .SP(clk_in_c_enable_58), .CK(clk_in_c), 
            .Q(s_7_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_7_2_c.GSR = "ENABLED";
    FD1P3AX s_7_3_c (.D(n645), .SP(clk_in_c_enable_58), .CK(clk_in_c), 
            .Q(s_7_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_7_3_c.GSR = "ENABLED";
    FD1P3AX s_7_4_c (.D(n649), .SP(clk_in_c_enable_58), .CK(clk_in_c), 
            .Q(s_7_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_7_4_c.GSR = "ENABLED";
    FD1P3AX s_7_5_c (.D(n653), .SP(clk_in_c_enable_58), .CK(clk_in_c), 
            .Q(s_7_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_7_5_c.GSR = "ENABLED";
    FD1P3AX s_7_6_c (.D(n657), .SP(clk_in_c_enable_58), .CK(clk_in_c), 
            .Q(s_7_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_7_6_c.GSR = "ENABLED";
    FD1S3AX s_7_7_c (.D(n661), .CK(clk_in_c), .Q(s_7_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_7_7_c.GSR = "ENABLED";
    FD1S3AX s_8_0_c (.D(n665), .CK(clk_in_c), .Q(s_8_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_8_0_c.GSR = "ENABLED";
    FD1P3AX s_8_1_c (.D(n669), .SP(clk_in_c_enable_64), .CK(clk_in_c), 
            .Q(s_8_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_8_1_c.GSR = "ENABLED";
    FD1P3AX s_8_2_c (.D(n673), .SP(clk_in_c_enable_64), .CK(clk_in_c), 
            .Q(s_8_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_8_2_c.GSR = "ENABLED";
    FD1P3AX s_8_3_c (.D(n677), .SP(clk_in_c_enable_64), .CK(clk_in_c), 
            .Q(s_8_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_8_3_c.GSR = "ENABLED";
    FD1P3AX s_8_4_c (.D(n681), .SP(clk_in_c_enable_64), .CK(clk_in_c), 
            .Q(s_8_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_8_4_c.GSR = "ENABLED";
    FD1P3AX s_8_5_c (.D(n685), .SP(clk_in_c_enable_64), .CK(clk_in_c), 
            .Q(s_8_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_8_5_c.GSR = "ENABLED";
    FD1P3AX s_8_6_c (.D(n689), .SP(clk_in_c_enable_64), .CK(clk_in_c), 
            .Q(s_8_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_8_6_c.GSR = "ENABLED";
    FD1S3AX s_8_7_c (.D(n693), .CK(clk_in_c), .Q(s_8_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_8_7_c.GSR = "ENABLED";
    FD1S3AX s_9_0_c (.D(n697), .CK(clk_in_c), .Q(s_9_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_9_0_c.GSR = "ENABLED";
    FD1P3AX s_9_1_c (.D(n701), .SP(clk_in_c_enable_70), .CK(clk_in_c), 
            .Q(s_9_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_9_1_c.GSR = "ENABLED";
    FD1P3AX s_9_2_c (.D(n714), .SP(clk_in_c_enable_70), .CK(clk_in_c), 
            .Q(s_9_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_9_2_c.GSR = "ENABLED";
    FD1P3AX s_9_3_c (.D(n718), .SP(clk_in_c_enable_70), .CK(clk_in_c), 
            .Q(s_9_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_9_3_c.GSR = "ENABLED";
    FD1P3AX s_9_4_c (.D(n722), .SP(clk_in_c_enable_70), .CK(clk_in_c), 
            .Q(s_9_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_9_4_c.GSR = "ENABLED";
    FD1P3AX s_9_5_c (.D(n726), .SP(clk_in_c_enable_70), .CK(clk_in_c), 
            .Q(s_9_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_9_5_c.GSR = "ENABLED";
    FD1P3AX s_9_6_c (.D(n730), .SP(clk_in_c_enable_70), .CK(clk_in_c), 
            .Q(s_9_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_9_6_c.GSR = "ENABLED";
    FD1S3AX s_9_7_c (.D(n734), .CK(clk_in_c), .Q(s_9_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_9_7_c.GSR = "ENABLED";
    FD1S3AX s_10_0_c (.D(n738), .CK(clk_in_c), .Q(s_10_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_10_0_c.GSR = "ENABLED";
    FD1P3AX s_10_1_c (.D(n742), .SP(clk_in_c_enable_76), .CK(clk_in_c), 
            .Q(s_10_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_10_1_c.GSR = "ENABLED";
    FD1P3AX s_10_2_c (.D(n746), .SP(clk_in_c_enable_76), .CK(clk_in_c), 
            .Q(s_10_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_10_2_c.GSR = "ENABLED";
    FD1P3AX s_10_3_c (.D(n750), .SP(clk_in_c_enable_76), .CK(clk_in_c), 
            .Q(s_10_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_10_3_c.GSR = "ENABLED";
    FD1P3AX s_10_4_c (.D(n754), .SP(clk_in_c_enable_76), .CK(clk_in_c), 
            .Q(s_10_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_10_4_c.GSR = "ENABLED";
    FD1P3AX s_10_5_c (.D(n758), .SP(clk_in_c_enable_76), .CK(clk_in_c), 
            .Q(s_10_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_10_5_c.GSR = "ENABLED";
    FD1P3AX s_10_6_c (.D(n762), .SP(clk_in_c_enable_76), .CK(clk_in_c), 
            .Q(s_10_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_10_6_c.GSR = "ENABLED";
    FD1S3AX s_10_7_c (.D(n766), .CK(clk_in_c), .Q(s_10_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_10_7_c.GSR = "ENABLED";
    FD1S3AX s_11_0_c (.D(n770), .CK(clk_in_c), .Q(s_11_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_11_0_c.GSR = "ENABLED";
    FD1P3AX s_11_1_c (.D(n774), .SP(clk_in_c_enable_82), .CK(clk_in_c), 
            .Q(s_11_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_11_1_c.GSR = "ENABLED";
    FD1P3AX s_11_2_c (.D(n778), .SP(clk_in_c_enable_82), .CK(clk_in_c), 
            .Q(s_11_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_11_2_c.GSR = "ENABLED";
    FD1P3AX s_11_3_c (.D(n782), .SP(clk_in_c_enable_82), .CK(clk_in_c), 
            .Q(s_11_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_11_3_c.GSR = "ENABLED";
    FD1P3AX s_11_4_c (.D(n786), .SP(clk_in_c_enable_82), .CK(clk_in_c), 
            .Q(s_11_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_11_4_c.GSR = "ENABLED";
    FD1P3AX s_11_5_c (.D(n790), .SP(clk_in_c_enable_82), .CK(clk_in_c), 
            .Q(s_11_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_11_5_c.GSR = "ENABLED";
    FD1P3AX s_11_6_c (.D(n794), .SP(clk_in_c_enable_82), .CK(clk_in_c), 
            .Q(s_11_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_11_6_c.GSR = "ENABLED";
    FD1S3AX s_11_7_c (.D(n798), .CK(clk_in_c), .Q(s_11_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_11_7_c.GSR = "ENABLED";
    FD1S3AX s_12_0_c (.D(n802), .CK(clk_in_c), .Q(s_12_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_12_0_c.GSR = "ENABLED";
    FD1P3AX s_12_1_c (.D(n806), .SP(clk_in_c_enable_88), .CK(clk_in_c), 
            .Q(s_12_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_12_1_c.GSR = "ENABLED";
    FD1P3AX s_12_2_c (.D(n810), .SP(clk_in_c_enable_88), .CK(clk_in_c), 
            .Q(s_12_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_12_2_c.GSR = "ENABLED";
    FD1P3AX s_12_3_c (.D(n814), .SP(clk_in_c_enable_88), .CK(clk_in_c), 
            .Q(s_12_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_12_3_c.GSR = "ENABLED";
    FD1P3AX s_12_4_c (.D(n818), .SP(clk_in_c_enable_88), .CK(clk_in_c), 
            .Q(s_12_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_12_4_c.GSR = "ENABLED";
    FD1P3AX s_12_5_c (.D(n822), .SP(clk_in_c_enable_88), .CK(clk_in_c), 
            .Q(s_12_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_12_5_c.GSR = "ENABLED";
    FD1P3AX s_12_6_c (.D(n826), .SP(clk_in_c_enable_88), .CK(clk_in_c), 
            .Q(s_12_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_12_6_c.GSR = "ENABLED";
    FD1S3AX s_12_7_c (.D(n830), .CK(clk_in_c), .Q(s_12_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_12_7_c.GSR = "ENABLED";
    FD1S3AX s_13_0_c (.D(n834), .CK(clk_in_c), .Q(s_13_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_13_0_c.GSR = "ENABLED";
    FD1P3AX s_13_1_c (.D(n838), .SP(clk_in_c_enable_94), .CK(clk_in_c), 
            .Q(s_13_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_13_1_c.GSR = "ENABLED";
    FD1P3AX s_13_2_c (.D(n842), .SP(clk_in_c_enable_94), .CK(clk_in_c), 
            .Q(s_13_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_13_2_c.GSR = "ENABLED";
    FD1P3AX s_13_3_c (.D(n846), .SP(clk_in_c_enable_94), .CK(clk_in_c), 
            .Q(s_13_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_13_3_c.GSR = "ENABLED";
    FD1P3AX s_13_4_c (.D(n850), .SP(clk_in_c_enable_94), .CK(clk_in_c), 
            .Q(s_13_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_13_4_c.GSR = "ENABLED";
    FD1P3AX s_13_5_c (.D(n854), .SP(clk_in_c_enable_94), .CK(clk_in_c), 
            .Q(s_13_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_13_5_c.GSR = "ENABLED";
    FD1P3AX s_13_6_c (.D(n858), .SP(clk_in_c_enable_94), .CK(clk_in_c), 
            .Q(s_13_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_13_6_c.GSR = "ENABLED";
    FD1S3AX s_13_7_c (.D(n862), .CK(clk_in_c), .Q(s_13_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_13_7_c.GSR = "ENABLED";
    FD1S3AX s_14_0_c (.D(n866), .CK(clk_in_c), .Q(s_14_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_14_0_c.GSR = "ENABLED";
    FD1P3AX s_14_1_c (.D(n870), .SP(clk_in_c_enable_100), .CK(clk_in_c), 
            .Q(s_14_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_14_1_c.GSR = "ENABLED";
    FD1P3AX s_14_2_c (.D(n874), .SP(clk_in_c_enable_100), .CK(clk_in_c), 
            .Q(s_14_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_14_2_c.GSR = "ENABLED";
    FD1P3AX s_14_3_c (.D(n878), .SP(clk_in_c_enable_100), .CK(clk_in_c), 
            .Q(s_14_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_14_3_c.GSR = "ENABLED";
    FD1P3AX s_14_4_c (.D(n882), .SP(clk_in_c_enable_100), .CK(clk_in_c), 
            .Q(s_14_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_14_4_c.GSR = "ENABLED";
    FD1P3AX s_14_5_c (.D(n886), .SP(clk_in_c_enable_100), .CK(clk_in_c), 
            .Q(s_14_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_14_5_c.GSR = "ENABLED";
    FD1P3AX s_14_6_c (.D(n890), .SP(clk_in_c_enable_100), .CK(clk_in_c), 
            .Q(s_14_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_14_6_c.GSR = "ENABLED";
    FD1S3AX s_14_7_c (.D(n894), .CK(clk_in_c), .Q(s_14_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_14_7_c.GSR = "ENABLED";
    FD1S3AX s_15_0_c (.D(n898), .CK(clk_in_c), .Q(s_15_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_15_0_c.GSR = "ENABLED";
    FD1P3AX s_15_1_c (.D(n902), .SP(clk_in_c_enable_106), .CK(clk_in_c), 
            .Q(s_15_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_15_1_c.GSR = "ENABLED";
    FD1P3AX s_15_2_c (.D(n906), .SP(clk_in_c_enable_106), .CK(clk_in_c), 
            .Q(s_15_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_15_2_c.GSR = "ENABLED";
    FD1P3AX s_15_3_c (.D(n910), .SP(clk_in_c_enable_106), .CK(clk_in_c), 
            .Q(s_15_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_15_3_c.GSR = "ENABLED";
    FD1P3AX s_15_4_c (.D(n914), .SP(clk_in_c_enable_106), .CK(clk_in_c), 
            .Q(s_15_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_15_4_c.GSR = "ENABLED";
    FD1P3AX s_15_5_c (.D(n918), .SP(clk_in_c_enable_106), .CK(clk_in_c), 
            .Q(s_15_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_15_5_c.GSR = "ENABLED";
    FD1P3AX s_15_6_c (.D(n922), .SP(clk_in_c_enable_106), .CK(clk_in_c), 
            .Q(s_15_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_15_6_c.GSR = "ENABLED";
    FD1S3AX s_15_7_c (.D(n926), .CK(clk_in_c), .Q(s_15_7)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam s_15_7_c.GSR = "ENABLED";
    FD1S3AX stack_1018 (.D(n1844[5]), .CK(clk_in_c), .Q(n2335));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1018.GSR = "ENABLED";
    PFUMX PrioSelect_473_i19 (.BLUT(n15_adj_474), .ALUT(n17_adj_475), .C0(n18993), 
          .Z(n814)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16531 (.D0(n19699), .D1(n19700), .SD(instruction[10]), .Z(n7_adj_476));
    PFUMX PrioSelect_469_i19 (.BLUT(n15_adj_477), .ALUT(n17_adj_478), .C0(n18993), 
          .Z(n810)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    CCU2D add_632_3 (.A0(instruction[1]), .B0(n7_adj_479), .C0(instruction[11]), 
          .D0(n14_adj_480), .A1(instruction[2]), .B1(n7_adj_481), .C1(instruction[11]), 
          .D1(n14_adj_482), .CIN(n14261), .COUT(n14262), .S0(Z_N_367[1]), 
          .S1(Z_N_367[2]));   // f:/home/mini-mcu/step_fpga/mcu.v(263[59:70])
    defparam add_632_3.INIT0 = 16'h56a6;
    defparam add_632_3.INIT1 = 16'h56a6;
    defparam add_632_3.INJECT1_0 = "NO";
    defparam add_632_3.INJECT1_1 = "NO";
    PFUMX PrioSelect_465_i19 (.BLUT(n15_adj_483), .ALUT(n17_adj_484), .C0(n18993), 
          .Z(n806)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1S1I out_port_7__I_0_i3 (.D(s_N_294[2]), .CK(out_port_7__N_232), .CD(n10012), 
           .Q(out_port[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam out_port_7__I_0_i3.GSR = "ENABLED";
    FD1S1I out_port_7__I_0_i4 (.D(s_N_294[3]), .CK(out_port_7__N_232), .CD(n10012), 
           .Q(out_port[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam out_port_7__I_0_i4.GSR = "ENABLED";
    FD1S1I out_port_7__I_0_i5 (.D(s_N_294[4]), .CK(out_port_7__N_232), .CD(n10012), 
           .Q(out_port[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam out_port_7__I_0_i5.GSR = "ENABLED";
    FD1S1I out_port_7__I_0_i6 (.D(s_N_294[5]), .CK(out_port_7__N_232), .CD(n10012), 
           .Q(out_port[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam out_port_7__I_0_i6.GSR = "ENABLED";
    FD1S1I out_port_7__I_0_i7 (.D(s_N_294[6]), .CK(out_port_7__N_232), .CD(n10012), 
           .Q(out_port[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam out_port_7__I_0_i7.GSR = "ENABLED";
    FD1S1I out_port_7__I_0_i8 (.D(C_N_336[0]), .CK(out_port_7__N_232), .CD(n10012), 
           .Q(out_port[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam out_port_7__I_0_i8.GSR = "ENABLED";
    FD1S1I port_id_7__I_0_i2 (.D(n23), .CK(port_id_7__N_215), .CD(n10010), 
           .Q(port_id[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam port_id_7__I_0_i2.GSR = "ENABLED";
    FD1S1I port_id_7__I_0_i3 (.D(n23_adj_485), .CK(port_id_7__N_215), .CD(n10010), 
           .Q(port_id[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam port_id_7__I_0_i3.GSR = "ENABLED";
    FD1S1I port_id_7__I_0_i4 (.D(n23_adj_486), .CK(port_id_7__N_215), .CD(n10010), 
           .Q(port_id[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam port_id_7__I_0_i4.GSR = "ENABLED";
    FD1S1I port_id_7__I_0_i5 (.D(n23_adj_487), .CK(port_id_7__N_215), .CD(n10010), 
           .Q(port_id[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam port_id_7__I_0_i5.GSR = "ENABLED";
    FD1S1I port_id_7__I_0_i6 (.D(n23_adj_488), .CK(port_id_7__N_215), .CD(n10010), 
           .Q(port_id[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam port_id_7__I_0_i6.GSR = "ENABLED";
    FD1S1I port_id_7__I_0_i7 (.D(n23_adj_489), .CK(port_id_7__N_215), .CD(n10010), 
           .Q(port_id[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam port_id_7__I_0_i7.GSR = "ENABLED";
    FD1S1I port_id_7__I_0_i8 (.D(n23_adj_490), .CK(port_id_7__N_215), .CD(n10010), 
           .Q(port_id[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam port_id_7__I_0_i8.GSR = "ENABLED";
    FD1S3AX stack_1017 (.D(n1844[4]), .CK(clk_in_c), .Q(n2333));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1017.GSR = "ENABLED";
    PFUMX PrioSelect_457_i16 (.BLUT(n14_adj_491), .ALUT(n15_adj_492), .C0(n18838), 
          .Z(n16_adj_493)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1S3AX stack_1016 (.D(n1844[3]), .CK(clk_in_c), .Q(n2331));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1016.GSR = "ENABLED";
    LUT4 i17338_3_lut_4_lut (.A(n22219), .B(n22102), .C(n14_adj_494), 
         .D(n10_c), .Z(n15_adj_495)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17338_3_lut_4_lut.init = 16'hf1e0;
    PFUMX PrioSelect_457_i13 (.BLUT(n8_adj_496), .ALUT(n12), .C0(n18826), 
          .Z(n13_adj_497)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_453_i19 (.BLUT(n15_adj_498), .ALUT(n17_adj_499), .C0(n18809), 
          .Z(n794)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1S3AX stack_1014 (.D(n1844[1]), .CK(clk_in_c), .Q(n2327));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1014.GSR = "ENABLED";
    FD1P3IX write_strobe_501 (.D(write_strobe_N_287), .SP(clk_in_c_enable_109), 
            .CD(n2730), .CK(clk_in_c), .Q(write_strobe));   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam write_strobe_501.GSR = "ENABLED";
    CCU2D add_632_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(instruction[0]), .B1(n7_adj_500), .C1(instruction[11]), 
          .D1(n14_adj_501), .COUT(n14261), .S1(Z_N_367[0]));   // f:/home/mini-mcu/step_fpga/mcu.v(263[59:70])
    defparam add_632_1.INIT0 = 16'hF000;
    defparam add_632_1.INIT1 = 16'h56a6;
    defparam add_632_1.INJECT1_0 = "NO";
    defparam add_632_1.INJECT1_1 = "NO";
    CCU2D add_21_5 (.A0(address[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(address[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14266), .COUT(n14267), .S0(n18[3]), .S1(n18[4]));   // f:/home/mini-mcu/step_fpga/mcu.v(217[27:35])
    defparam add_21_5.INIT0 = 16'h5aaa;
    defparam add_21_5.INIT1 = 16'h5aaa;
    defparam add_21_5.INJECT1_0 = "NO";
    defparam add_21_5.INJECT1_1 = "NO";
    PFUMX PrioSelect_449_i19 (.BLUT(n15_adj_502), .ALUT(n17_adj_503), .C0(n18809), 
          .Z(n790)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_445_i19 (.BLUT(n15_adj_504), .ALUT(n17_adj_505), .C0(n18809), 
          .Z(n786)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_441_i19 (.BLUT(n15_adj_506), .ALUT(n17_adj_507), .C0(n18809), 
          .Z(n782)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17751_4_lut (.A(n22151), .B(n22153), .C(n22152), .D(n213[4]), 
         .Z(n17550)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17751_4_lut.init = 16'haaab;
    FD1S3AX stack_1013 (.D(n1844[0]), .CK(clk_in_c), .Q(n2325));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1013.GSR = "ENABLED";
    PFUMX PrioSelect_437_i19 (.BLUT(n15_adj_508), .ALUT(n17_adj_509), .C0(n18809), 
          .Z(n778)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1S3AX stack_1015 (.D(n1844[2]), .CK(clk_in_c), .Q(n2329));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1015.GSR = "ENABLED";
    PFUMX PrioSelect_433_i19 (.BLUT(n15_adj_510), .ALUT(n17_adj_511), .C0(n18809), 
          .Z(n774)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1P3AX i123_124 (.D(C), .SP(n1[20]), .CK(clk_in_c), .Q(stack_zc_d0_20_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i123_124.GSR = "ENABLED";
    PFUMX PrioSelect_425_i16 (.BLUT(n14_adj_512), .ALUT(n15_adj_513), .C0(n18654), 
          .Z(n16_adj_514)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i3226_3_lut_4_lut (.A(n22227), .B(n22281), .C(n13_adj_515), .D(n13_adj_516), 
         .Z(n10_adj_517)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i3226_3_lut_4_lut.init = 16'hf780;
    FD1S3AX stack_1012 (.D(clk_in_c_enable_115), .CK(clk_in_c), .Q(n2322));   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam stack_1012.GSR = "ENABLED";
    FD1P3IX enable_intr_flag_507 (.D(instruction[0]), .SP(clk_in_c_enable_113), 
            .CD(n22301), .CK(clk_in_c), .Q(enable_intr_flag));   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam enable_intr_flag_507.GSR = "ENABLED";
    SPR16X4C creg0 (.DI0(s_N_294[4]), .DI1(s_N_294[5]), .DI2(s_N_294[6]), 
            .DI3(C_N_336[0]), .AD0(instruction[0]), .AD1(instruction[1]), 
            .AD2(instruction[2]), .AD3(instruction[3]), .CK(clk_in_c), 
            .WRE(creg_N_407), .DO0(n1108[4]), .DO1(n1108[5]), .DO2(n1108[6]), 
            .DO3(n1108[7]));
    defparam creg0.initval = "0x0000000000000000";
    FD1S3AX stack_1010 (.D(n3[4]), .CK(clk_in_c), .Q(n2320));   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam stack_1010.GSR = "ENABLED";
    FD1P3AX i117_118 (.D(C), .SP(n1[19]), .CK(clk_in_c), .Q(stack_zc_d0_19_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i117_118.GSR = "ENABLED";
    LUT4 PrioSelect_181_i11_3_lut_4_lut (.A(n22235), .B(n11714), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_519)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_181_i11_3_lut_4_lut.init = 16'hfd20;
    FD1S3AX stack (.D(n1844[11]), .CK(clk_in_c), .Q(n2347));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack.GSR = "ENABLED";
    PDPW8KC stack0 (.DI0(n1844[0]), .DI1(n1844[1]), .DI2(n1844[2]), .DI3(n1844[3]), 
            .DI4(n1844[4]), .DI5(n1844[5]), .DI6(n1844[6]), .DI7(n1844[7]), 
            .DI8(n1844[8]), .DI9(n1844[9]), .DI10(n1844[10]), .DI11(n1844[11]), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(stack_N_397[0]), .ADW1(stack_N_397[1]), 
            .ADW2(stack_N_397[2]), .ADW3(n22288), .ADW4(stack_N_397[4]), 
            .ADW5(GND_net), .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), 
            .BE0(VCC_net), .BE1(VCC_net), .CEW(clk_in_c_enable_115), .CLKW(clk_in_c), 
            .CSW0(GND_net), .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), 
            .ADR1(GND_net), .ADR2(GND_net), .ADR3(GND_net), .ADR4(n3[0]), 
            .ADR5(n3[1]), .ADR6(n3[2]), .ADR7(n3[3]), .ADR8(n3[4]), 
            .ADR9(GND_net), .ADR10(GND_net), .ADR11(GND_net), .ADR12(GND_net), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(clk_in_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n2342), 
            .DO1(n2344), .DO2(n2346), .DO9(n2324), .DO10(n2326), .DO11(n2328), 
            .DO12(n2330), .DO13(n2332), .DO14(n2334), .DO15(n2336), 
            .DO16(n2338), .DO17(n2340));
    defparam stack0.DATA_WIDTH_W = 18;
    defparam stack0.DATA_WIDTH_R = 18;
    defparam stack0.REGMODE = "NOREG";
    defparam stack0.CSDECODE_W = "0b000";
    defparam stack0.CSDECODE_R = "0b000";
    defparam stack0.GSR = "DISABLED";
    defparam stack0.RESETMODE = "SYNC";
    defparam stack0.ASYNC_RESET_RELEASE = "SYNC";
    defparam stack0.INIT_DATA = "STATIC";
    defparam stack0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam stack0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    LUT4 PrioSelect_245_i13_3_lut_4_lut (.A(n22259), .B(n7762), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_520)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_245_i13_3_lut_4_lut.init = 16'hf780;
    FD1S3AX stack_1023 (.D(n1844[10]), .CK(clk_in_c), .Q(n2345));   // f:/home/mini-mcu/step_fpga/mcu.v(284[36:45])
    defparam stack_1023.GSR = "ENABLED";
    FD1P3AX i111_112 (.D(C), .SP(n1[18]), .CK(clk_in_c), .Q(stack_zc_d0_18_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i111_112.GSR = "ENABLED";
    FD1P3AX i105_106 (.D(C), .SP(n1[17]), .CK(clk_in_c), .Q(stack_zc_d0_17_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i105_106.GSR = "ENABLED";
    FD1P3AX i99_100 (.D(C), .SP(n1[16]), .CK(clk_in_c), .Q(stack_zc_d0_16_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i99_100.GSR = "ENABLED";
    PFUMX PrioSelect_421_i19 (.BLUT(n15_adj_521), .ALUT(n17_adj_522), .C0(n18625), 
          .Z(n762)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_417_i19 (.BLUT(n15_adj_523), .ALUT(n17_adj_524), .C0(n18625), 
          .Z(n758)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1P3AX i93_94 (.D(C), .SP(n1[15]), .CK(clk_in_c), .Q(stack_zc_d0_15_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i93_94.GSR = "ENABLED";
    FD1P3AX i87_88 (.D(C), .SP(n1[14]), .CK(clk_in_c), .Q(stack_zc_d0_14_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i87_88.GSR = "ENABLED";
    FD1P3AX i81_82 (.D(C), .SP(n1[13]), .CK(clk_in_c), .Q(stack_zc_d0_13_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i81_82.GSR = "ENABLED";
    FD1P3AX i75_76 (.D(C), .SP(n1[12]), .CK(clk_in_c), .Q(stack_zc_d0_12_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i75_76.GSR = "ENABLED";
    FD1P3AX i69_70 (.D(C), .SP(n1[11]), .CK(clk_in_c), .Q(stack_zc_d0_11_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i69_70.GSR = "ENABLED";
    FD1P3AX i63_64 (.D(C), .SP(n1[10]), .CK(clk_in_c), .Q(stack_zc_d0_10_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i63_64.GSR = "ENABLED";
    FD1P3AX i57_58 (.D(C), .SP(n1[9]), .CK(clk_in_c), .Q(stack_zc_d0_9_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i57_58.GSR = "ENABLED";
    FD1P3AX i51_52 (.D(C), .SP(n1[8]), .CK(clk_in_c), .Q(stack_zc_d0_8_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i51_52.GSR = "ENABLED";
    FD1P3AX i45_46 (.D(C), .SP(n1[7]), .CK(clk_in_c), .Q(stack_zc_d0_7_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i45_46.GSR = "ENABLED";
    FD1P3AX i39_40 (.D(C), .SP(n1[6]), .CK(clk_in_c), .Q(stack_zc_d0_6_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i39_40.GSR = "ENABLED";
    FD1P3AX i33_34 (.D(C), .SP(n1[5]), .CK(clk_in_c), .Q(stack_zc_d0_5_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i33_34.GSR = "ENABLED";
    PFUMX PrioSelect_413_i19 (.BLUT(n15_adj_525), .ALUT(n17_adj_526), .C0(n18625), 
          .Z(n754)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1P3AX i27_28 (.D(C), .SP(n1[4]), .CK(clk_in_c), .Q(stack_zc_d0_4_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i27_28.GSR = "ENABLED";
    FD1P3AX i21_22 (.D(C), .SP(n1[3]), .CK(clk_in_c), .Q(stack_zc_d0_3_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i21_22.GSR = "ENABLED";
    FD1P3AX i15_16 (.D(C), .SP(n1[2]), .CK(clk_in_c), .Q(stack_zc_d0_2_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i15_16.GSR = "ENABLED";
    FD1P3AX i9_10 (.D(C), .SP(n1[1]), .CK(clk_in_c), .Q(stack_zc_d0_1_0));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i9_10.GSR = "ENABLED";
    FD1P3AX i126_127 (.D(Z), .SP(n1[20]), .CK(clk_in_c), .Q(stack_zc_20_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i126_127.GSR = "ENABLED";
    LUT4 PrioSelect_497_i12_3_lut_4_lut (.A(n22254), .B(n7908), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_527)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_497_i12_3_lut_4_lut.init = 16'hf780;
    FD1P3AX i120_121 (.D(Z), .SP(n1[19]), .CK(clk_in_c), .Q(stack_zc_19_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i120_121.GSR = "ENABLED";
    FD1P3AX i114_115 (.D(Z), .SP(n1[18]), .CK(clk_in_c), .Q(stack_zc_18_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i114_115.GSR = "ENABLED";
    FD1P3AX i108_109 (.D(Z), .SP(n1[17]), .CK(clk_in_c), .Q(stack_zc_17_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i108_109.GSR = "ENABLED";
    FD1P3AX i102_103 (.D(Z), .SP(n1[16]), .CK(clk_in_c), .Q(stack_zc_16_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i102_103.GSR = "ENABLED";
    LUT4 i17336_3_lut_4_lut (.A(n22219), .B(n22102), .C(n14_adj_528), 
         .D(n10_adj_529), .Z(n15_adj_530)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17336_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX i96_97 (.D(Z), .SP(n1[15]), .CK(clk_in_c), .Q(stack_zc_15_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i96_97.GSR = "ENABLED";
    FD1P3AX i90_91 (.D(Z), .SP(n1[14]), .CK(clk_in_c), .Q(stack_zc_14_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i90_91.GSR = "ENABLED";
    LUT4 PrioSelect_85_i14_3_lut_4_lut_4_lut (.A(n11714), .B(n13_adj_531), 
         .C(Z_N_387[2]), .D(n22251), .Z(n14_adj_532)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_85_i14_3_lut_4_lut_4_lut.init = 16'hccd8;
    FD1P3AX i84_85 (.D(Z), .SP(n1[13]), .CK(clk_in_c), .Q(stack_zc_13_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i84_85.GSR = "ENABLED";
    LUT4 PrioSelect_77_i5_3_lut_4_lut (.A(n8627), .B(n11714), .C(n7_adj_479), 
         .D(n7_adj_473), .Z(n5)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_77_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17769_4_lut (.A(n22151), .B(n22153), .C(n22152), .D(n17508), 
         .Z(n20371)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17769_4_lut.init = 16'habaa;
    FD1P3AX i78_79 (.D(Z), .SP(n1[12]), .CK(clk_in_c), .Q(stack_zc_12_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i78_79.GSR = "ENABLED";
    FD1P3AX i72_73 (.D(Z), .SP(n1[11]), .CK(clk_in_c), .Q(stack_zc_11_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i72_73.GSR = "ENABLED";
    FD1P3AX i66_67 (.D(Z), .SP(n1[10]), .CK(clk_in_c), .Q(stack_zc_10_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i66_67.GSR = "ENABLED";
    FD1P3AX i60_61 (.D(Z), .SP(n1[9]), .CK(clk_in_c), .Q(stack_zc_9_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i60_61.GSR = "ENABLED";
    FD1P3AX i54_55 (.D(Z), .SP(n1[8]), .CK(clk_in_c), .Q(stack_zc_8_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i54_55.GSR = "ENABLED";
    PFUMX PrioSelect_409_i19 (.BLUT(n15_adj_533), .ALUT(n17_adj_534), .C0(n18625), 
          .Z(n750)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1P3AX i48_49 (.D(Z), .SP(n1[7]), .CK(clk_in_c), .Q(stack_zc_7_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i48_49.GSR = "ENABLED";
    FD1P3AX i42_43 (.D(Z), .SP(n1[6]), .CK(clk_in_c), .Q(stack_zc_6_1));   // f:/home/mini-mcu/step_fpga/mcu.v(118[44:52])
    defparam i42_43.GSR = "ENABLED";
    PFUMX PrioSelect_405_i19 (.BLUT(n15_adj_535), .ALUT(n17_adj_536), .C0(n18625), 
          .Z(n746)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i14318_4_lut (.A(n22150), .B(n22149), .C(n22148), .D(n213[4]), 
         .Z(n17508)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14318_4_lut.init = 16'h5554;
    PFUMX PrioSelect_401_i19 (.BLUT(n15_adj_537), .ALUT(n17_adj_538), .C0(n18625), 
          .Z(n742)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_1_lut_rep_732 (.A(jp), .Z(n22299)) /* synthesis lut_function=(!(A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_1_lut_rep_732.init = 16'h5555;
    PFUMX PrioSelect_393_i16 (.BLUT(n14_adj_539), .ALUT(n15_adj_540), .C0(n18321), 
          .Z(n16_adj_541)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_501_i12_3_lut_4_lut (.A(n22254), .B(n7908), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_542)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_501_i12_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_393_i13 (.BLUT(n8_adj_543), .ALUT(n12_adj_544), .C0(n18306), 
          .Z(n13_adj_545)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1S3AX st__i1 (.D(n3[1]), .CK(clk_in_c), .Q(st[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam st__i1.GSR = "ENABLED";
    L6MUX21 i16538 (.D0(n19706), .D1(n19707), .SD(instruction[10]), .Z(n7_adj_473));
    PFUMX PrioSelect_389_i19 (.BLUT(n15_adj_546), .ALUT(n17_adj_547), .C0(n18361), 
          .Z(n730)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    CCU2D add_412_3 (.A0(instruction[1]), .B0(instruction[11]), .C0(n7_adj_479), 
          .D0(n14_adj_480), .A1(instruction[2]), .B1(instruction[11]), 
          .C1(n7_adj_481), .D1(n14_adj_482), .CIN(n14274), .COUT(n14275), 
          .S0(Z_N_378[1]), .S1(Z_N_378[2]));   // f:/home/mini-mcu/step_fpga/mcu.v(275[74:85])
    defparam add_412_3.INIT0 = 16'ha965;
    defparam add_412_3.INIT1 = 16'ha965;
    defparam add_412_3.INJECT1_0 = "NO";
    defparam add_412_3.INJECT1_1 = "NO";
    PFUMX PrioSelect_385_i19 (.BLUT(n15_adj_548), .ALUT(n17_adj_549), .C0(n18361), 
          .Z(n726)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_381_i19 (.BLUT(n15_adj_550), .ALUT(n17_adj_551), .C0(n18361), 
          .Z(n722)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_377_i19 (.BLUT(n15_adj_552), .ALUT(n17_adj_553), .C0(n18361), 
          .Z(n718)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    CCU2D add_827_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14286), 
          .S0(C_N_342[8]));   // f:/home/mini-mcu/step_fpga/mcu.v(281[97:106])
    defparam add_827_cout.INIT0 = 16'h0000;
    defparam add_827_cout.INIT1 = 16'h0000;
    defparam add_827_cout.INJECT1_0 = "NO";
    defparam add_827_cout.INJECT1_1 = "NO";
    CCU2D add_412_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(instruction[0]), .B1(instruction[11]), .C1(n7_adj_500), 
          .D1(n14_adj_501), .COUT(n14274), .S1(Z_N_378[0]));   // f:/home/mini-mcu/step_fpga/mcu.v(275[74:85])
    defparam add_412_1.INIT0 = 16'h0000;
    defparam add_412_1.INIT1 = 16'ha965;
    defparam add_412_1.INJECT1_0 = "NO";
    defparam add_412_1.INJECT1_1 = "NO";
    PFUMX PrioSelect_373_i19 (.BLUT(n15_adj_554), .ALUT(n17_adj_555), .C0(n18361), 
          .Z(n714)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_369_i19 (.BLUT(n15_adj_556), .ALUT(n17_adj_557), .C0(n18361), 
          .Z(n701)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1S3AX st__i2 (.D(n3[2]), .CK(clk_in_c), .Q(st[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam st__i2.GSR = "ENABLED";
    FD1S3AX st__i3 (.D(n3[3]), .CK(clk_in_c), .Q(st[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam st__i3.GSR = "ENABLED";
    FD1S3AX st__i4 (.D(n3[4]), .CK(clk_in_c), .Q(st[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam st__i4.GSR = "ENABLED";
    FD1S3IX intr_f__i1 (.D(intr_f[0]), .CK(clk_in_c), .CD(n22301), .Q(intr_f[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(154[8] 157[4])
    defparam intr_f__i1.GSR = "ENABLED";
    FD1S3IX intr_f__i2 (.D(intr_f[1]), .CK(clk_in_c), .CD(n22301), .Q(intr_f[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(154[8] 157[4])
    defparam intr_f__i2.GSR = "ENABLED";
    FD1P3IX st_zc__i1 (.D(n2755), .SP(clk_in_c_enable_159), .CD(n22301), 
            .CK(clk_in_c), .Q(st_zc[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam st_zc__i1.GSR = "ENABLED";
    PFUMX PrioSelect_361_i16 (.BLUT(n14_adj_558), .ALUT(n15_adj_559), .C0(n18286), 
          .Z(n16_adj_560)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_357_i19 (.BLUT(n15_adj_561), .ALUT(n17_adj_562), .C0(n18257), 
          .Z(n689)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1P3IX st_zc__i2 (.D(n2634[1]), .SP(clk_in_c_enable_159), .CD(n22301), 
            .CK(clk_in_c), .Q(st_zc[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam st_zc__i2.GSR = "ENABLED";
    FD1P3IX st_zc__i3 (.D(n22316), .SP(clk_in_c_enable_159), .CD(n22301), 
            .CK(clk_in_c), .Q(st_zc[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam st_zc__i3.GSR = "ENABLED";
    FD1P3IX st_zc__i4 (.D(n2634[3]), .SP(clk_in_c_enable_159), .CD(n22301), 
            .CK(clk_in_c), .Q(st_zc[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam st_zc__i4.GSR = "ENABLED";
    LUT4 PrioSelect_505_i12_3_lut_4_lut (.A(n22254), .B(n7908), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_563)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_505_i12_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_353_i19 (.BLUT(n15_adj_564), .ALUT(n17_adj_565), .C0(n18257), 
          .Z(n685)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_349_i19 (.BLUT(n15_adj_566), .ALUT(n17_adj_567), .C0(n18257), 
          .Z(n681)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_345_i19 (.BLUT(n15_adj_568), .ALUT(n17_adj_569), .C0(n18257), 
          .Z(n677)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1P3IX pc__i2 (.D(n1238[1]), .SP(clk_in_c_enable_175), .CD(n10021), 
            .CK(clk_in_c), .Q(address[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i2.GSR = "ENABLED";
    PFUMX PrioSelect_341_i19 (.BLUT(n15_adj_570), .ALUT(n17_adj_571), .C0(n18257), 
          .Z(n673)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_337_i19 (.BLUT(n15_adj_572), .ALUT(n17_adj_573), .C0(n18257), 
          .Z(n669)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1P3JX pc__i3 (.D(n1238[2]), .SP(clk_in_c_enable_175), .PD(n10021), 
            .CK(clk_in_c), .Q(address[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i3.GSR = "ENABLED";
    FD1P3IX pc__i4 (.D(n1238[3]), .SP(clk_in_c_enable_175), .CD(n10021), 
            .CK(clk_in_c), .Q(address[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i4.GSR = "ENABLED";
    PFUMX PrioSelect_329_i16 (.BLUT(n14_adj_574), .ALUT(n15_adj_575), .C0(n18102), 
          .Z(n16_adj_576)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1P3JX pc__i5 (.D(n1238[4]), .SP(clk_in_c_enable_175), .PD(n10021), 
            .CK(clk_in_c), .Q(address[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i5.GSR = "ENABLED";
    FD1P3IX pc__i6 (.D(n1238[5]), .SP(clk_in_c_enable_175), .CD(n10021), 
            .CK(clk_in_c), .Q(address[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i6.GSR = "ENABLED";
    FD1P3JX pc__i7 (.D(n1238[6]), .SP(clk_in_c_enable_175), .PD(n10021), 
            .CK(clk_in_c), .Q(address[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i7.GSR = "ENABLED";
    PFUMX PrioSelect_329_i13 (.BLUT(n8_adj_577), .ALUT(n12_adj_578), .C0(n18090), 
          .Z(n13_adj_579)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1P3IX pc__i8 (.D(n1238[7]), .SP(clk_in_c_enable_175), .CD(n10021), 
            .CK(clk_in_c), .Q(address[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i8.GSR = "ENABLED";
    FD1P3IX pc__i9 (.D(n1238[8]), .SP(clk_in_c_enable_175), .CD(n10021), 
            .CK(clk_in_c), .Q(address[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i9.GSR = "ENABLED";
    FD1P3IX pc__i10 (.D(n1238[9]), .SP(clk_in_c_enable_175), .CD(n10021), 
            .CK(clk_in_c), .Q(address[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i10.GSR = "ENABLED";
    FD1P3IX pc__i11 (.D(n1238[10]), .SP(clk_in_c_enable_175), .CD(n10021), 
            .CK(clk_in_c), .Q(address[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i11.GSR = "ENABLED";
    LUT4 PrioSelect_509_i12_3_lut_4_lut (.A(n22254), .B(n7908), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_580)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_509_i12_3_lut_4_lut.init = 16'hf780;
    FD1P3IX pc__i12 (.D(n1238[11]), .SP(clk_in_c_enable_175), .CD(n10021), 
            .CK(clk_in_c), .Q(address[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i12.GSR = "ENABLED";
    FD1P3IX pc__i13 (.D(n18[12]), .SP(clk_in_c_enable_175), .CD(n21516), 
            .CK(clk_in_c), .Q(pc[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i13.GSR = "ENABLED";
    PFUMX PrioSelect_325_i19 (.BLUT(n15_adj_581), .ALUT(n17_adj_582), .C0(n18073), 
          .Z(n657)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_513_i12_3_lut_4_lut (.A(n22254), .B(n7908), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_583)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_513_i12_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_321_i19 (.BLUT(n15_adj_584), .ALUT(n17_adj_585), .C0(n18073), 
          .Z(n653)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17640_2_lut_rep_562_3_lut_4_lut_4_lut (.A(n11714), .B(n11778), 
         .C(n22277), .D(n10_adj_586), .Z(n22129)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i17640_2_lut_rep_562_3_lut_4_lut_4_lut.init = 16'h0001;
    PFUMX PrioSelect_317_i19 (.BLUT(n15_adj_587), .ALUT(n17_adj_588), .C0(n18073), 
          .Z(n649)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_313_i19 (.BLUT(n15_adj_589), .ALUT(n17_adj_590), .C0(n18073), 
          .Z(n645)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_309_i19 (.BLUT(n15_adj_591), .ALUT(n17_adj_592), .C0(n18073), 
          .Z(n640)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    FD1P3IX C_506 (.D(C_N_304), .SP(clk_in_c_enable_173), .CD(n22301), 
            .CK(clk_in_c), .Q(C));   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam C_506.GSR = "ENABLED";
    FD1S1I out_port_7__I_0_i2 (.D(s_N_294[1]), .CK(out_port_7__N_232), .CD(n10012), 
           .Q(out_port[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam out_port_7__I_0_i2.GSR = "ENABLED";
    FD1P3AX Z_509 (.D(Z_N_356), .SP(clk_in_c_enable_174), .CK(clk_in_c), 
            .Q(Z));   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam Z_509.GSR = "ENABLED";
    FD1S1I port_id_7__I_0_i1 (.D(n23_adj_593), .CK(port_id_7__N_215), .CD(n10010), 
           .Q(port_id[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam port_id_7__I_0_i1.GSR = "ENABLED";
    PFUMX PrioSelect_305_i19 (.BLUT(n15_adj_594), .ALUT(n17_adj_595), .C0(n18073), 
          .Z(n636)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1482_3_lut_4_lut (.A(n8627), .B(n11714), .C(n7_adj_481), .D(n7_adj_500), 
         .Z(n10_adj_596)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1482_3_lut_4_lut.init = 16'hfd20;
    FD1S1I out_port_7__I_0_i1 (.D(out_port_7__N_232), .CK(out_port_7__N_232), 
           .CD(n22228), .Q(out_port[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(403[1] 424[4])
    defparam out_port_7__I_0_i1.GSR = "ENABLED";
    FD1P3IX pc__i1 (.D(n1238[0]), .SP(clk_in_c_enable_175), .CD(n10021), 
            .CK(clk_in_c), .Q(address[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam pc__i1.GSR = "ENABLED";
    PFUMX PrioSelect_297_i16 (.BLUT(n14_adj_597), .ALUT(n15_adj_598), .C0(n17918), 
          .Z(n16_adj_599)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_293_i19 (.BLUT(n15_adj_600), .ALUT(n17_adj_601), .C0(n17889), 
          .Z(n624)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_269_i5_3_lut_4_lut (.A(n7762), .B(n8647), .C(n7_adj_479), 
         .D(n7_adj_473), .Z(n5_adj_602)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_269_i5_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_289_i19 (.BLUT(n15_adj_603), .ALUT(n17_adj_604), .C0(n17889), 
          .Z(n620)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_285_i19 (.BLUT(n15_adj_605), .ALUT(n17_adj_606), .C0(n17889), 
          .Z(n616)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_281_i19 (.BLUT(n15_adj_607), .ALUT(n17_adj_608), .C0(n17889), 
          .Z(n612)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16545 (.D0(n19713), .D1(n19714), .SD(instruction[10]), .Z(n7_adj_609));
    LUT4 i17474_4_lut (.A(n22145), .B(n22147), .C(n22146), .D(n213[3]), 
         .Z(n17366)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17474_4_lut.init = 16'haaab;
    PFUMX PrioSelect_277_i19 (.BLUT(n15_adj_610), .ALUT(n17_adj_611), .C0(n17889), 
          .Z(n608)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_273_i19 (.BLUT(n15_adj_612), .ALUT(n17_adj_613), .C0(n17889), 
          .Z(n604)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16552 (.D0(n19720), .D1(n19721), .SD(instruction[10]), .Z(n7_adj_462));
    PFUMX PrioSelect_265_i16 (.BLUT(n14_adj_614), .ALUT(n15_adj_615), .C0(n17734), 
          .Z(n16_adj_616)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i18407 (.BLUT(n22311), .ALUT(n22312), .C0(st[3]), .Z(n22313));
    PFUMX PrioSelect_265_i13 (.BLUT(n8_adj_617), .ALUT(n12_adj_618), .C0(n17722), 
          .Z(n13_adj_619)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_517_i12_3_lut_4_lut (.A(n22254), .B(n7908), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_620)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_517_i12_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_261_i19 (.BLUT(n15_adj_621), .ALUT(n17_adj_622), .C0(n17705), 
          .Z(n592)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_493_i15_3_lut_4_lut (.A(n22254), .B(n7908), .C(n1108[0]), 
         .D(n5_adj_623), .Z(n15_adj_624)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_493_i15_3_lut_4_lut.init = 16'hf780;
    L6MUX21 i16559 (.D0(n19727), .D1(n19728), .SD(instruction[10]), .Z(n7_c));
    LUT4 PrioSelect_89_i14_3_lut_4_lut_4_lut (.A(n11714), .B(n13_adj_625), 
         .C(Z_N_387[3]), .D(n22251), .Z(n14_adj_626)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_89_i14_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX PrioSelect_257_i19 (.BLUT(n15_adj_627), .ALUT(n17_adj_628), .C0(n17705), 
          .Z(n588)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_253_i19 (.BLUT(n15_adj_629), .ALUT(n17_adj_630), .C0(n17705), 
          .Z(n575)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_521_i15_3_lut_4_lut (.A(n22254), .B(n7908), .C(n1108[7]), 
         .D(n9_adj_631), .Z(n15_adj_632)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_521_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i8439_4_lut (.A(s_3_7), .B(n16278), .C(n7_adj_476), .D(n16246), 
         .Z(n6)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8439_4_lut.init = 16'h3022;
    PFUMX PrioSelect_249_i19 (.BLUT(n15_adj_633), .ALUT(n17_adj_634), .C0(n17705), 
          .Z(n571)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_245_i19 (.BLUT(n15_adj_635), .ALUT(n17_adj_636), .C0(n17705), 
          .Z(n567)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16566 (.D0(n19734), .D1(n19735), .SD(instruction[10]), .Z(n7_adj_500));
    PFUMX PrioSelect_241_i19 (.BLUT(n15_adj_637), .ALUT(n17_adj_638), .C0(n17705), 
          .Z(n563)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_233_i16 (.BLUT(n14_adj_639), .ALUT(n15_adj_640), .C0(n17550), 
          .Z(n16_adj_641)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_229_i19 (.BLUT(n15_adj_642), .ALUT(n17_adj_643), .C0(n17521), 
          .Z(n551)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_225_i19 (.BLUT(n15_adj_644), .ALUT(n17_adj_645), .C0(n17521), 
          .Z(n547)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_221_i19 (.BLUT(n15_adj_646), .ALUT(n17_adj_647), .C0(n17521), 
          .Z(n543)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_77_i14_3_lut_4_lut_4_lut (.A(n11714), .B(n10_adj_648), 
         .C(Z_N_387[0]), .D(n22251), .Z(n14_adj_649)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_77_i14_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX PrioSelect_217_i19 (.BLUT(n15_adj_650), .ALUT(n17_adj_651), .C0(n17521), 
          .Z(n539)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_105_i14_3_lut_4_lut_4_lut (.A(n11714), .B(n10_adj_652), 
         .C(Z_N_387[7]), .D(n22251), .Z(n14_adj_653)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_105_i14_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_177_i11_3_lut_4_lut (.A(n22235), .B(n11714), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_654)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_177_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_93_i14_3_lut_4_lut_4_lut (.A(n11714), .B(n13_adj_655), 
         .C(Z_N_387[4]), .D(n22251), .Z(n14_adj_656)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_93_i14_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_81_i14_3_lut_4_lut_4_lut (.A(n11714), .B(n13_adj_657), 
         .C(Z_N_387[1]), .D(n22251), .Z(n14_adj_658)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_81_i14_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_97_i14_3_lut_4_lut_4_lut (.A(n11714), .B(n13_adj_659), 
         .C(Z_N_387[5]), .D(n22251), .Z(n14_adj_660)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_97_i14_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_101_i14_3_lut_4_lut_4_lut (.A(n11714), .B(n13_adj_661), 
         .C(Z_N_387[6]), .D(n22251), .Z(n14_adj_662)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_101_i14_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_185_i11_3_lut_4_lut (.A(n22235), .B(n11714), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_663)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_185_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_189_i11_3_lut_4_lut (.A(n22235), .B(n11714), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_664)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_189_i11_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_213_i19 (.BLUT(n15_adj_665), .ALUT(n17_adj_666), .C0(n17521), 
          .Z(n535)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_209_i19 (.BLUT(n15_adj_667), .ALUT(n17_adj_668), .C0(n17521), 
          .Z(n531)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_201_i16 (.BLUT(n14_adj_669), .ALUT(n15_adj_670), .C0(n17366), 
          .Z(n16_adj_671)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_193_i11_3_lut_4_lut (.A(n22235), .B(n11714), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_672)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_193_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_197_i11_3_lut_4_lut (.A(n22235), .B(n11714), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_673)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_197_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17529_4_lut (.A(n22145), .B(n22147), .C(n22146), .D(n17324), 
         .Z(n20131)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17529_4_lut.init = 16'habaa;
    PFUMX PrioSelect_201_i13 (.BLUT(n8_c), .ALUT(n12_adj_674), .C0(n17354), 
          .Z(n13_adj_675)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_197_i19 (.BLUT(n15_adj_676), .ALUT(n17_adj_677), .C0(n17337), 
          .Z(n519)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i14134_4_lut (.A(n22144), .B(n22143), .C(n22142), .D(n213[3]), 
         .Z(n17324)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14134_4_lut.init = 16'h5554;
    LUT4 PrioSelect_501_i11_3_lut_4_lut (.A(n22255), .B(n7908), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_678)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_501_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_193_i19 (.BLUT(n15_adj_679), .ALUT(n17_adj_680), .C0(n17337), 
          .Z(n515)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_497_i11_3_lut_4_lut (.A(n22255), .B(n7908), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_681)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_497_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_505_i11_3_lut_4_lut (.A(n22255), .B(n7908), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_682)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_505_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i17579_4_lut (.A(n22139), .B(n22141), .C(n22140), .D(n213[2]), 
         .Z(n17182)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17579_4_lut.init = 16'haaab;
    PFUMX PrioSelect_189_i19 (.BLUT(n15_adj_683), .ALUT(n17_adj_684), .C0(n17337), 
          .Z(n511)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_509_i11_3_lut_4_lut (.A(n22255), .B(n7908), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_685)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_509_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_513_i11_3_lut_4_lut (.A(n22255), .B(n7908), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_686)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_513_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_517_i11_3_lut_4_lut (.A(n22255), .B(n7908), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_687)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_517_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut (.A(st_zc[1]), .B(n22284), .C(n7746), .D(n22307), 
         .Z(n1[17])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 PrioSelect_201_i11_3_lut_4_lut (.A(n22236), .B(n11714), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_688)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_201_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17597_4_lut (.A(n22139), .B(n22141), .C(n22140), .D(n17140), 
         .Z(n20199)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17597_4_lut.init = 16'habaa;
    L6MUX21 i18220 (.D0(n21794), .D1(n21791), .SD(instruction[1]), .Z(n21795));
    LUT4 i13950_4_lut (.A(n22138), .B(n22137), .C(n22136), .D(n213[2]), 
         .Z(n17140)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i13950_4_lut.init = 16'h5554;
    LUT4 i1_2_lut_3_lut_4_lut_adj_34 (.A(st_zc[1]), .B(n22284), .C(n22285), 
         .D(n22307), .Z(n1[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_34.init = 16'h0400;
    PFUMX i18218 (.BLUT(n21793), .ALUT(n21792), .C0(instruction[3]), .Z(n21794));
    LUT4 i1_2_lut_3_lut_4_lut_adj_35 (.A(st_zc[1]), .B(n22284), .C(n22282), 
         .D(n22307), .Z(n1[13])) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_35.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_36 (.A(st_zc[1]), .B(n22284), .C(n22285), 
         .D(n22307), .Z(n1[1])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_36.init = 16'h0004;
    LUT4 PrioSelect_493_i11_3_lut_4_lut (.A(n22253), .B(n7908), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_689)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_493_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_185_i19 (.BLUT(n15_adj_690), .ALUT(n17_adj_691), .C0(n17337), 
          .Z(n507)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_adj_37 (.A(st_zc[1]), .B(n22284), .C(n22282), 
         .D(n22307), .Z(n1[9])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_37.init = 16'h0040;
    LUT4 PrioSelect_521_i11_3_lut_4_lut (.A(n22253), .B(n7908), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_692)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_521_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_550_3_lut_4_lut (.A(n7908), .B(n7876), .C(n16417), 
         .D(n160), .Z(n22117)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_rep_550_3_lut_4_lut.init = 16'h8000;
    LUT4 PrioSelect_173_i11_3_lut_4_lut (.A(n22236), .B(n11714), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_693)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_173_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17699_4_lut (.A(n22133), .B(n22135), .C(n22134), .D(n213[1]), 
         .Z(n16998)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17699_4_lut.init = 16'haaab;
    LUT4 i1_2_lut_3_lut_4_lut_adj_38 (.A(n22304), .B(n22283), .C(n22282), 
         .D(n22307), .Z(n1[8])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_38.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_39 (.A(n22304), .B(n22283), .C(n22285), 
         .D(n22307), .Z(n1[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_39.init = 16'h0400;
    PFUMX i18214 (.BLUT(n21790), .ALUT(n21789), .C0(instruction[3]), .Z(n21791));
    LUT4 i8421_4_lut (.A(s_1_7), .B(n16279), .C(n7_adj_476), .D(n16251), 
         .Z(n6_adj_694)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8421_4_lut.init = 16'h3022;
    LUT4 i1_2_lut_3_lut_4_lut_adj_40 (.A(n22304), .B(n22283), .C(n22282), 
         .D(n22307), .Z(n1[12])) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_40.init = 16'h4000;
    LUT4 i16784_3_lut (.A(stack_zc_14_1), .B(stack_zc_15_1), .C(st_zc[0]), 
         .Z(n19954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16784_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_697_3_lut_3_lut_4_lut (.A(clk_in_c_enable_174), .B(instruction[15]), 
         .C(n8070), .D(n8_adj_695), .Z(n22264)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_697_3_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i16783_3_lut (.A(stack_zc_12_1), .B(stack_zc_13_1), .C(st_zc[0]), 
         .Z(n19953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16783_3_lut.init = 16'hcaca;
    LUT4 i16782_3_lut (.A(stack_zc_10_1), .B(stack_zc_11_1), .C(st_zc[0]), 
         .Z(n19952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16782_3_lut.init = 16'hcaca;
    LUT4 i16781_3_lut (.A(stack_zc_8_1), .B(stack_zc_9_1), .C(st_zc[0]), 
         .Z(n19951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16781_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_241_i13_3_lut_4_lut (.A(n22259), .B(n7762), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_696)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_241_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_660_4_lut (.A(n206), .B(instruction[0]), .C(instruction[3]), 
         .D(n7646), .Z(n22227)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i1_2_lut_rep_660_4_lut.init = 16'hb000;
    LUT4 PrioSelect_241_i14_3_lut_4_lut (.A(n22257), .B(n7762), .C(Z_N_387[1]), 
         .D(n13_adj_696), .Z(n14_adj_697)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_241_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i13421_2_lut_rep_699_3_lut_3_lut_4_lut (.A(clk_in_c_enable_174), 
         .B(instruction[14]), .C(instruction[13]), .D(n10_adj_698), .Z(n22266)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i13421_2_lut_rep_699_3_lut_3_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_3_lut (.A(instruction[1]), .B(instruction[2]), .C(instruction[0]), 
         .Z(n160)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i1_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i16780_3_lut (.A(stack_zc_6_1), .B(stack_zc_7_1), .C(st_zc[0]), 
         .Z(n19950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16780_3_lut.init = 16'hcaca;
    LUT4 i16779_3_lut (.A(stack_zc_4_1), .B(stack_zc_5_1), .C(st_zc[0]), 
         .Z(n19949)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16779_3_lut.init = 16'hcaca;
    LUT4 i2378_3_lut_4_lut (.A(n8627), .B(n16312), .C(n14_adj_482), .D(n14_adj_501), 
         .Z(n10_adj_699)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2378_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_245_i14_3_lut_4_lut (.A(n22257), .B(n7762), .C(Z_N_387[2]), 
         .D(n13_adj_520), .Z(n14_adj_700)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_245_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i2394_3_lut_4_lut (.A(n8627), .B(n16312), .C(n14), .D(n14_adj_480), 
         .Z(n10_adj_701)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2394_3_lut_4_lut.init = 16'hf780;
    LUT4 i2410_3_lut_4_lut (.A(n8627), .B(n16312), .C(n14_adj_463), .D(n14_adj_482), 
         .Z(n10_adj_702)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2410_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_249_i14_3_lut_4_lut (.A(n22257), .B(n7762), .C(Z_N_387[3]), 
         .D(n13_adj_703), .Z(n14_adj_704)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_249_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i16778_3_lut (.A(stack_zc_2_1), .B(stack_zc_3_1), .C(st_zc[0]), 
         .Z(n19948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16778_3_lut.init = 16'hcaca;
    LUT4 i16777_3_lut (.A(stack_zc_1_1), .B(st_zc[0]), .Z(n19947)) /* synthesis lut_function=(A (B)) */ ;
    defparam i16777_3_lut.init = 16'h8888;
    LUT4 i16769_3_lut (.A(stack_zc_d0_14_0), .B(stack_zc_d0_15_0), .C(st_zc[0]), 
         .Z(n19939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16769_3_lut.init = 16'hcaca;
    LUT4 i16768_3_lut (.A(stack_zc_d0_12_0), .B(stack_zc_d0_13_0), .C(st_zc[0]), 
         .Z(n19938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16768_3_lut.init = 16'hcaca;
    LUT4 i2426_3_lut_4_lut (.A(n8627), .B(n16312), .C(n14_adj_705), .D(n14), 
         .Z(n10_adj_706)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2426_3_lut_4_lut.init = 16'hf780;
    LUT4 i8842_2_lut_rep_696_3_lut_3_lut_4_lut (.A(clk_in_c_enable_174), .B(instruction[15]), 
         .C(n9_adj_707), .D(n8_adj_708), .Z(n22263)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i8842_2_lut_rep_696_3_lut_3_lut_4_lut.init = 16'hfffd;
    LUT4 i2442_3_lut_4_lut (.A(n8627), .B(n16312), .C(n14_adj_709), .D(n14_adj_463), 
         .Z(n10_adj_710)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2442_3_lut_4_lut.init = 16'hf780;
    LUT4 i16767_3_lut (.A(stack_zc_d0_10_0), .B(stack_zc_d0_11_0), .C(st_zc[0]), 
         .Z(n19937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16767_3_lut.init = 16'hcaca;
    LUT4 i2458_3_lut_4_lut (.A(n8627), .B(n16312), .C(n14_adj_711), .D(n14_adj_705), 
         .Z(n10_adj_712)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2458_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_397_i5_3_lut_4_lut (.A(n8647), .B(n16312), .C(n14_adj_480), 
         .D(n14_adj_711), .Z(n5_adj_713)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_397_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i16766_3_lut (.A(stack_zc_d0_8_0), .B(stack_zc_d0_9_0), .C(st_zc[0]), 
         .Z(n19936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16766_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_253_i14_3_lut_4_lut (.A(n22257), .B(n7762), .C(Z_N_387[4]), 
         .D(n13_adj_714), .Z(n14_adj_715)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_253_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i16765_3_lut (.A(stack_zc_d0_6_0), .B(stack_zc_d0_7_0), .C(st_zc[0]), 
         .Z(n19935)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16765_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_4_lut (.A(s_N_294[1]), .B(instruction[1]), .C(s_N_294[2]), 
         .D(instruction[2]), .Z(n10_adj_716)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(429[15:76])
    defparam i2_2_lut_4_lut.init = 16'h7888;
    LUT4 PrioSelect_257_i14_3_lut_4_lut (.A(n22257), .B(n7762), .C(Z_N_387[5]), 
         .D(n13_adj_717), .Z(n14_adj_718)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_257_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i16764_3_lut (.A(stack_zc_d0_4_0), .B(stack_zc_d0_5_0), .C(st_zc[0]), 
         .Z(n19934)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16764_3_lut.init = 16'hcaca;
    LUT4 i2602_3_lut_4_lut (.A(n8647), .B(n16312), .C(n14_adj_482), .D(n14_adj_501), 
         .Z(n10_adj_719)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2602_3_lut_4_lut.init = 16'hf780;
    LUT4 i16763_3_lut (.A(stack_zc_d0_2_0), .B(stack_zc_d0_3_0), .C(st_zc[0]), 
         .Z(n19933)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16763_3_lut.init = 16'hcaca;
    LUT4 i16762_3_lut (.A(stack_zc_d0_1_0), .B(st_zc[0]), .Z(n19932)) /* synthesis lut_function=(A (B)) */ ;
    defparam i16762_3_lut.init = 16'h8888;
    LUT4 i17658_2_lut_rep_522_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n16392), 
         .C(n7762), .D(n22268), .Z(n22089)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17658_2_lut_rep_522_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i16760_3_lut (.A(stack_zc_d0_18_0), .B(stack_zc_d0_19_0), .C(st_zc[0]), 
         .Z(n19930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16760_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_41 (.A(instruction[10]), .B(instruction[11]), 
         .C(instruction[9]), .Z(n8044)) /* synthesis lut_function=(A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_3_lut_adj_41.init = 16'h8080;
    LUT4 i16759_3_lut (.A(stack_zc_d0_16_0), .B(stack_zc_d0_17_0), .C(st_zc[0]), 
         .Z(n19929)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16759_3_lut.init = 16'hcaca;
    LUT4 i2618_3_lut_4_lut (.A(n8647), .B(n16312), .C(n14), .D(n14_adj_480), 
         .Z(n10_adj_720)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2618_3_lut_4_lut.init = 16'hf780;
    LUT4 i16757_3_lut (.A(stack_zc_18_1), .B(stack_zc_19_1), .C(st_zc[0]), 
         .Z(n19927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16757_3_lut.init = 16'hcaca;
    LUT4 i16756_3_lut (.A(stack_zc_16_1), .B(stack_zc_17_1), .C(st_zc[0]), 
         .Z(n19926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16756_3_lut.init = 16'hcaca;
    LUT4 n2083_bdd_4_lut_17852 (.A(n22109), .B(n2085), .C(n16312), .D(n11778), 
         .Z(n21081)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;
    defparam n2083_bdd_4_lut_17852.init = 16'hff1f;
    LUT4 PrioSelect_521_i8_4_lut (.A(n6_adj_721), .B(n14_adj_711), .C(n7925), 
         .D(n7921), .Z(n8_adj_722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_521_i8_4_lut.init = 16'hcfca;
    PFUMX PrioSelect_181_i19 (.BLUT(n15_adj_723), .ALUT(n17_adj_724), .C0(n17337), 
          .Z(n503)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17766_2_lut_rep_527_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n16392), 
         .C(n16312), .D(n22268), .Z(n22094)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17766_2_lut_rep_527_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 PrioSelect_261_i14_3_lut_4_lut (.A(n22257), .B(n7762), .C(Z_N_387[6]), 
         .D(n13_adj_725), .Z(n14_adj_726)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_261_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17594_2_lut_rep_532_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n16392), 
         .C(n7908), .D(n22268), .Z(n22099)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17594_2_lut_rep_532_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i2634_3_lut_4_lut (.A(n8647), .B(n16312), .C(n14_adj_463), .D(n14_adj_482), 
         .Z(n10_adj_727)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2634_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_714_4_lut (.A(instruction[10]), .B(instruction[11]), 
         .C(instruction[8]), .D(instruction[9]), .Z(n22281)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_rep_714_4_lut.init = 16'h8000;
    LUT4 i2650_3_lut_4_lut (.A(n8647), .B(n16312), .C(n14_adj_705), .D(n14), 
         .Z(n10_adj_728)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2650_3_lut_4_lut.init = 16'hf780;
    LUT4 i2666_3_lut_4_lut (.A(n8647), .B(n16312), .C(n14_adj_709), .D(n14_adj_463), 
         .Z(n10_adj_729)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2666_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_42 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n7762), .Z(n54[7])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_42.init = 16'h8000;
    LUT4 i2682_3_lut_4_lut (.A(n8647), .B(n16312), .C(n14_adj_711), .D(n14_adj_705), 
         .Z(n10_adj_730)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2682_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_461_i5_3_lut_4_lut (.A(n8627), .B(n7908), .C(n13_adj_731), 
         .D(n14_adj_711), .Z(n5_adj_732)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_461_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_237_i14_3_lut_4_lut (.A(n22257), .B(n7762), .C(Z_N_387[0]), 
         .D(n10_adj_733), .Z(n14_adj_734)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_237_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_265_i14_3_lut_4_lut (.A(n22257), .B(n7762), .C(Z_N_387[7]), 
         .D(n10_adj_735), .Z(n14_adj_614)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_265_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_43 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n16312), .Z(n16349)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_43.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_44 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n7908), .Z(n7946)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_44.init = 16'h8000;
    LUT4 i2826_3_lut_4_lut (.A(n8627), .B(n7908), .C(n13_adj_736), .D(n5_adj_737), 
         .Z(n10_adj_738)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2826_3_lut_4_lut.init = 16'hf780;
    LUT4 i2842_3_lut_4_lut (.A(n8627), .B(n7908), .C(n13_adj_739), .D(n13_adj_731), 
         .Z(n10_adj_740)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2842_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_45 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n11714), .Z(n16258)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_45.init = 16'h0080;
    LUT4 i2858_3_lut_4_lut (.A(n8627), .B(n7908), .C(n13_adj_516), .D(n13_adj_736), 
         .Z(n10_adj_741)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2858_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_46 (.A(n2071), .B(instruction[9]), .C(instruction[8]), 
         .D(n16312), .Z(n16355)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_46.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_47 (.A(n2071), .B(instruction[9]), .C(instruction[8]), 
         .D(n7908), .Z(n7945)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_47.init = 16'h0800;
    PFUMX PrioSelect_177_i19 (.BLUT(n15_adj_742), .ALUT(n17_adj_743), .C0(n17337), 
          .Z(n499)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_adj_48 (.A(n2071), .B(instruction[9]), .C(instruction[8]), 
         .D(n7762), .Z(n54[6])) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_48.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_49 (.A(n2071), .B(instruction[9]), .C(instruction[8]), 
         .D(n11714), .Z(n16244)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_49.init = 16'h0008;
    LUT4 i2874_3_lut_4_lut (.A(n8627), .B(n7908), .C(n13_adj_744), .D(n13_adj_739), 
         .Z(n10_adj_745)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2874_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_50 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n7908), .Z(n7944)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_50.init = 16'h0800;
    LUT4 PrioSelect_277_i11_3_lut_4_lut (.A(n22229), .B(n7762), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_746)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_277_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_51 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n11714), .Z(n16259)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_51.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_52 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n16312), .Z(n16350)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_52.init = 16'h0800;
    LUT4 i2890_3_lut_4_lut (.A(n8627), .B(n7908), .C(n13_adj_515), .D(n13_adj_516), 
         .Z(n10_adj_747)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2890_3_lut_4_lut.init = 16'hf780;
    LUT4 i2906_3_lut_4_lut (.A(n8627), .B(n7908), .C(n13_adj_748), .D(n13_adj_744), 
         .Z(n10_adj_749)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2906_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_53 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n7762), .Z(n54[5])) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_53.init = 16'h0800;
    LUT4 i17540_2_lut_2_lut_3_lut_4_lut_3_lut_4_lut (.A(instruction[11]), 
         .B(instruction[10]), .C(n22246), .D(n22250), .Z(n16727)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;
    defparam i17540_2_lut_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h0111;
    LUT4 i1_2_lut_3_lut_4_lut_adj_54 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n7762), .Z(n151[4])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_54.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_55 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n16312), .Z(n16341)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_55.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_56 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n11714), .Z(n16268)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_56.init = 16'h0002;
    LUT4 PrioSelect_105_i9_3_lut_4_lut (.A(n22101), .B(n11714), .C(n7_adj_500), 
         .D(C), .Z(n9_c)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_105_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13350_2_lut_4_lut (.A(s_N_294[4]), .B(instruction[4]), .C(s_N_294[5]), 
         .D(instruction[5]), .Z(n16508)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;
    defparam i13350_2_lut_4_lut.init = 16'hf888;
    LUT4 i17182_3_lut_4_lut (.A(n22135), .B(n22084), .C(n14_adj_750), 
         .D(n10_adj_751), .Z(n15_adj_752)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17182_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i121_4_lut_3_lut (.A(instruction[13]), .B(instruction[14]), .C(instruction[15]), 
         .Z(n55)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i121_4_lut_3_lut.init = 16'h4242;
    LUT4 PrioSelect_273_i11_3_lut_4_lut (.A(n22229), .B(n7762), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_753)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_273_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i13371_2_lut_4_lut (.A(C_N_336[0]), .B(instruction[7]), .C(out_port_7__N_217[0]), 
         .D(instruction[0]), .Z(n16532)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;
    defparam i13371_2_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut (.A(instruction[17]), .B(instruction[16]), .C(instruction[14]), 
         .D(instruction[13]), .Z(n66)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_3_lut_4_lut.init = 16'haaa8;
    PFUMX PrioSelect_169_i16 (.BLUT(n14_adj_754), .ALUT(n15_adj_755), .C0(n17182), 
          .Z(n16_adj_756)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17172_3_lut_4_lut (.A(n22135), .B(n22084), .C(n14_adj_757), 
         .D(n10_adj_758), .Z(n15_adj_759)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17172_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17178_3_lut_4_lut (.A(n22135), .B(n22084), .C(n14_adj_760), 
         .D(n10_adj_761), .Z(n15_adj_762)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17178_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_281_i11_3_lut_4_lut (.A(n22229), .B(n7762), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_763)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_281_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_3_lut_4_lut (.A(instruction[16]), .B(instruction[14]), .C(instruction[13]), 
         .D(n56), .Z(n14413)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_57 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n7908), .Z(n7926)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_57.init = 16'h0200;
    LUT4 PrioSelect_285_i11_3_lut_4_lut (.A(n22229), .B(n7762), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_764)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_285_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_289_i11_3_lut_4_lut (.A(n22229), .B(n7762), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_765)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_289_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_293_i11_3_lut_4_lut (.A(n22229), .B(n7762), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_766)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_293_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_58 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n7908), .Z(n7943)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_58.init = 16'h0200;
    LUT4 instruction_17__I_0_568_i11_2_lut_rep_712_4_lut (.A(instruction[12]), 
         .B(n8050), .C(instruction[15]), .D(n9_adj_707), .Z(n22279)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[17:23])
    defparam instruction_17__I_0_568_i11_2_lut_rep_712_4_lut.init = 16'hffdf;
    LUT4 i17176_3_lut_4_lut (.A(n22135), .B(n22084), .C(n14_adj_767), 
         .D(n10_adj_768), .Z(n15_adj_769)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17176_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17180_3_lut_4_lut (.A(n22135), .B(n22084), .C(n14_adj_770), 
         .D(n10_adj_771), .Z(n15_adj_772)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17180_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17174_3_lut_4_lut (.A(n22135), .B(n22084), .C(n14_adj_773), 
         .D(n10_adj_774), .Z(n15_adj_775)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17174_3_lut_4_lut.init = 16'hf1e0;
    LUT4 instruction_17__I_0_557_i10_2_lut_3_lut (.A(instruction[15]), .B(instruction[16]), 
         .C(instruction[17]), .Z(n10_adj_776)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(240[16:24])
    defparam instruction_17__I_0_557_i10_2_lut_3_lut.init = 16'hefef;
    LUT4 PrioSelect_137_i9_3_lut_4_lut (.A(n22093), .B(n11714), .C(n7_adj_500), 
         .D(C), .Z(n9_adj_777)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_137_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17196_3_lut_4_lut (.A(n22141), .B(n22085), .C(n14_adj_778), 
         .D(n10_adj_779), .Z(n15_adj_780)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17196_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_59 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n11714), .Z(n16252)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_59.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_adj_60 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n16312), .Z(n16347)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_60.init = 16'h0200;
    LUT4 PrioSelect_553_i8_4_lut (.A(n6_adj_781), .B(n14_adj_711), .C(n7924), 
         .D(n7920), .Z(n8_adj_782)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_553_i8_4_lut.init = 16'hcfca;
    LUT4 i17186_3_lut_4_lut (.A(n22141), .B(n22085), .C(n14_adj_783), 
         .D(n10_adj_784), .Z(n15_adj_785)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17186_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17192_3_lut_4_lut (.A(n22141), .B(n22085), .C(n14_adj_786), 
         .D(n10_adj_787), .Z(n15_adj_788)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17192_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_61 (.A(n2071), .B(instruction[8]), .C(instruction[9]), 
         .D(n7762), .Z(n54[4])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(221[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_61.init = 16'h0200;
    LUT4 i17190_3_lut_4_lut (.A(n22141), .B(n22085), .C(n14_adj_790), 
         .D(n10_adj_791), .Z(n15_adj_792)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17190_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17194_3_lut_4_lut (.A(n22141), .B(n22085), .C(n14_adj_793), 
         .D(n10_adj_794), .Z(n15_adj_795)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17194_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_62 (.A(n2081), .B(instruction[9]), .C(instruction[8]), 
         .D(n11714), .Z(n16269)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_62.init = 16'h0008;
    LUT4 i1_2_lut (.A(instruction[10]), .B(instruction[11]), .Z(n7908)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_63 (.A(n2081), .B(instruction[9]), .C(instruction[8]), 
         .D(n16312), .Z(n16338)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_63.init = 16'h0800;
    PFUMX PrioSelect_165_i19 (.BLUT(n15_adj_780), .ALUT(n17_adj_796), .C0(n17153), 
          .Z(n487)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_adj_64 (.A(n2081), .B(instruction[9]), .C(instruction[8]), 
         .D(n7762), .Z(n151[6])) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_64.init = 16'h0800;
    LUT4 i17485_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22237), .B(n11714), .C(n22235), 
         .D(n22236), .Z(n17354)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17485_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3332;
    LUT4 i17188_3_lut_4_lut (.A(n22141), .B(n22085), .C(n14_adj_797), 
         .D(n10_adj_798), .Z(n15_adj_799)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17188_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n2083_bdd_4_lut_17857 (.A(n22109), .B(n2085), .C(n16312), .D(n7726), 
         .Z(n21098)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam n2083_bdd_4_lut_17857.init = 16'h1fff;
    LUT4 PrioSelect_169_i9_3_lut_4_lut (.A(n22095), .B(n11714), .C(n7_adj_500), 
         .D(C), .Z(n9_adj_800)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_169_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut_4_lut_adj_65 (.A(n2081), .B(instruction[9]), .C(instruction[8]), 
         .D(n7908), .Z(n7924)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_65.init = 16'h0800;
    LUT4 i17209_3_lut_4_lut (.A(n22147), .B(n22086), .C(n14_adj_801), 
         .D(n10_adj_802), .Z(n15_adj_676)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17209_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17199_3_lut_4_lut (.A(n22147), .B(n22086), .C(n14_adj_803), 
         .D(n10_adj_804), .Z(n15_adj_742)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17199_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17205_3_lut_4_lut (.A(n22147), .B(n22086), .C(n14_adj_805), 
         .D(n10_adj_806), .Z(n15_adj_683)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17205_3_lut_4_lut.init = 16'hf1e0;
    LUT4 instruction_17__I_0_569_i11_2_lut_rep_711_4_lut (.A(instruction[12]), 
         .B(n16484), .C(instruction[15]), .D(n9_adj_707), .Z(n22278)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[17:26])
    defparam instruction_17__I_0_569_i11_2_lut_rep_711_4_lut.init = 16'hffdf;
    LUT4 i17203_3_lut_4_lut (.A(n22147), .B(n22086), .C(n14_adj_807), 
         .D(n10_adj_808), .Z(n15_adj_690)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17203_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17207_3_lut_4_lut (.A(n22147), .B(n22086), .C(n14_adj_809), 
         .D(n10_adj_810), .Z(n15_adj_679)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17207_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_534_3_lut (.A(n2085), .B(instruction[8]), .C(instruction[9]), 
         .Z(n22101)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam i1_2_lut_rep_534_3_lut.init = 16'h0202;
    PFUMX PrioSelect_161_i19 (.BLUT(n15_adj_795), .ALUT(n17_adj_811), .C0(n17153), 
          .Z(n483)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_3_lut_4_lut_adj_66 (.A(clk_in_c_enable_109), .B(instruction[12]), 
         .C(n8050), .D(n10_adj_812), .Z(n4)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_3_lut_4_lut_adj_66.init = 16'haaa2;
    LUT4 i1_2_lut_rep_530_3_lut (.A(n2085), .B(instruction[8]), .C(instruction[9]), 
         .Z(n22097)) /* synthesis lut_function=(A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam i1_2_lut_rep_530_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_67 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n11714), .Z(n16283)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_67.init = 16'h0080;
    LUT4 instruction_17__I_0_555_i11_2_lut_rep_708_4_lut (.A(instruction[12]), 
         .B(n8050), .C(instruction[15]), .D(n8070), .Z(n22275)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(234[16:28])
    defparam instruction_17__I_0_555_i11_2_lut_rep_708_4_lut.init = 16'hfffe;
    PFUMX PrioSelect_157_i19 (.BLUT(n15_adj_788), .ALUT(n17_adj_813), .C0(n17153), 
          .Z(n479)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_173_i12_3_lut_4_lut (.A(n22237), .B(n11714), .C(Z_N_378[0]), 
         .D(n11_adj_693), .Z(n12_adj_814)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_173_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut_4_lut_adj_68 (.A(n22304), .B(n22283), .C(n7746), 
         .D(n22307), .Z(n1[16])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_68.init = 16'h0040;
    LUT4 i13482_4_lut_4_lut (.A(n22123), .B(n16644), .C(n22124), .D(n22125), 
         .Z(n16652)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i13482_4_lut_4_lut.init = 16'h0010;
    LUT4 n2083_bdd_4_lut_17821 (.A(n22109), .B(n2085), .C(n11714), .D(n7876), 
         .Z(n20976)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam n2083_bdd_4_lut_17821.init = 16'hf1ff;
    LUT4 i17779_3_lut_4_lut (.A(instruction[13]), .B(instruction[15]), .C(n9_adj_815), 
         .D(instruction[14]), .Z(write_strobe_N_287)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i17779_3_lut_4_lut.init = 16'h0400;
    PFUMX PrioSelect_153_i19 (.BLUT(n15_adj_792), .ALUT(n17_adj_816), .C0(n17153), 
          .Z(n475)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_adj_69 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n7908), .Z(n7923)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_69.init = 16'h8000;
    LUT4 i17201_3_lut_4_lut (.A(n22147), .B(n22086), .C(n14_adj_817), 
         .D(n10_adj_818), .Z(n15_adj_723)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17201_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_70 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n7762), .Z(n151[7])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_70.init = 16'h8000;
    LUT4 i17715_4_lut (.A(n22133), .B(n22135), .C(n22134), .D(n16956), 
         .Z(n20317)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17715_4_lut.init = 16'habaa;
    LUT4 i1_2_lut_3_lut_4_lut_adj_71 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n16312), .Z(n16331)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_71.init = 16'h8000;
    LUT4 PrioSelect_201_i9_3_lut_4_lut (.A(n22097), .B(n11714), .C(n7_adj_500), 
         .D(C), .Z(n9_adj_820)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_201_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17223_3_lut_4_lut (.A(n22153), .B(n22087), .C(n14_adj_821), 
         .D(n10_adj_822), .Z(n15_adj_642)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17223_3_lut_4_lut.init = 16'hf1e0;
    LUT4 instruction_17__I_0_556_i11_2_lut_rep_707_4_lut (.A(instruction[12]), 
         .B(n8050), .C(instruction[15]), .D(n8070), .Z(n22274)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[16:28])
    defparam instruction_17__I_0_556_i11_2_lut_rep_707_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_rep_706_4_lut (.A(instruction[12]), .B(n8050), .C(instruction[15]), 
         .D(n9_adj_707), .Z(n22273)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(216[16:21])
    defparam i1_2_lut_rep_706_4_lut.init = 16'hfffd;
    LUT4 instruction_17__I_0_530_i11_2_lut_rep_705_4_lut (.A(instruction[12]), 
         .B(n8050), .C(instruction[15]), .D(n8070), .Z(n22272)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(382[17:26])
    defparam instruction_17__I_0_530_i11_2_lut_rep_705_4_lut.init = 16'hffef;
    LUT4 i17213_3_lut_4_lut (.A(n22153), .B(n22087), .C(n14_adj_823), 
         .D(n10_adj_824), .Z(n15_adj_667)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17213_3_lut_4_lut.init = 16'hf1e0;
    PFUMX PrioSelect_149_i19 (.BLUT(n15_adj_799), .ALUT(n17_adj_825), .C0(n17153), 
          .Z(n471)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 instruction_17__I_0_553_i11_2_lut_rep_704_4_lut (.A(instruction[12]), 
         .B(n8050), .C(instruction[15]), .D(n8070), .Z(n22271)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(383[17:25])
    defparam instruction_17__I_0_553_i11_2_lut_rep_704_4_lut.init = 16'hffdf;
    LUT4 i1_2_lut_3_lut_adj_72 (.A(instruction[8]), .B(instruction[9]), 
         .C(n16378), .Z(clk_in_c_enable_58)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_72.init = 16'h8080;
    LUT4 i17219_3_lut_4_lut (.A(n22153), .B(n22087), .C(n14_adj_826), 
         .D(n10_adj_827), .Z(n15_adj_646)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17219_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_703_4_lut (.A(instruction[14]), .B(instruction[13]), 
         .C(instruction[15]), .D(n8070), .Z(n22270)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_703_4_lut.init = 16'hfffe;
    LUT4 PrioSelect_297_i11_3_lut_4_lut (.A(n22230), .B(n7762), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_828)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_297_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_528_3_lut (.A(n2085), .B(instruction[9]), .C(instruction[8]), 
         .Z(n22095)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam i1_2_lut_rep_528_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_3_lut_adj_73 (.A(instruction[8]), .B(instruction[9]), 
         .C(n16378), .Z(clk_in_c_enable_46)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_73.init = 16'h2020;
    LUT4 i13352_2_lut_rep_702_4_lut (.A(instruction[12]), .B(n8050), .C(instruction[16]), 
         .D(instruction[17]), .Z(n22269)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i13352_2_lut_rep_702_4_lut.init = 16'hffdf;
    LUT4 i13766_4_lut (.A(n22132), .B(n22131), .C(n22130), .D(n213[1]), 
         .Z(n16956)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i13766_4_lut.init = 16'h5554;
    LUT4 i2_3_lut_4_lut_adj_74 (.A(instruction[13]), .B(instruction[16]), 
         .C(Z), .D(Z_N_377), .Z(n14358)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i2_3_lut_4_lut_adj_74.init = 16'h8000;
    LUT4 i1_2_lut_rep_526_3_lut (.A(n2085), .B(instruction[8]), .C(instruction[9]), 
         .Z(n22093)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam i1_2_lut_rep_526_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_2_lut (.A(instruction[14]), .B(Z), .Z(n34)) /* synthesis lut_function=(!(A+!(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_75 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n11714), .Z(n16282)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_75.init = 16'h0008;
    PFUMX PrioSelect_145_i19 (.BLUT(n15_adj_785), .ALUT(n17_adj_829), .C0(n17153), 
          .Z(n467)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_adj_76 (.A(n22304), .B(n22283), .C(n7746), 
         .D(n22307), .Z(n1[20])) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_76.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_77 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n7908), .Z(n7925)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_77.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_78 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n16312), .Z(n16326)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_78.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_79 (.A(n2081), .B(instruction[8]), .C(instruction[9]), 
         .D(n7762), .Z(n151[5])) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(226[39:43])
    defparam i1_2_lut_3_lut_4_lut_adj_79.init = 16'h0800;
    LUT4 instruction_17__I_0_529_i10_2_lut_3_lut (.A(instruction[15]), .B(instruction[16]), 
         .C(instruction[17]), .Z(n10_adj_812)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(257[16:26])
    defparam instruction_17__I_0_529_i10_2_lut_3_lut.init = 16'hdfdf;
    LUT4 i1_3_lut_4_lut_adj_80 (.A(instruction[13]), .B(instruction[14]), 
         .C(instruction[12]), .D(n10_adj_812), .Z(n6978)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(363[17:25])
    defparam i1_3_lut_4_lut_adj_80.init = 16'hff7f;
    LUT4 i2_3_lut_4_lut_adj_81 (.A(instruction[13]), .B(instruction[14]), 
         .C(instruction[17]), .D(instruction[12]), .Z(n8_adj_830)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i2_3_lut_4_lut_adj_81.init = 16'h0004;
    LUT4 i17217_3_lut_4_lut (.A(n22153), .B(n22087), .C(n14_adj_831), 
         .D(n10_adj_832), .Z(n15_adj_650)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17217_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_655_3_lut_4_lut (.A(n160), .B(n7646), .C(instruction[11]), 
         .D(instruction[10]), .Z(n22222)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_655_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_82 (.A(n160), .B(n7646), .C(instruction[9]), 
         .D(instruction[8]), .Z(n15_adj_833)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_82.init = 16'h0080;
    LUT4 PrioSelect_269_i11_3_lut_4_lut (.A(n22230), .B(n7762), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_834)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_269_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut (.A(instruction[9]), .B(n8789), .C(instruction[11]), 
         .D(instruction[10]), .Z(n16253)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_4_lut.init = 16'h0004;
    LUT4 i17221_3_lut_4_lut (.A(n22153), .B(n22087), .C(n14_adj_835), 
         .D(n10_adj_836), .Z(n15_adj_644)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17221_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2_3_lut_3_lut (.A(instruction[16]), .B(instruction[14]), .C(C_N_338[8]), 
         .Z(n14422)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i2_3_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_4_lut_adj_83 (.A(instruction[9]), .B(n8789), .C(instruction[11]), 
         .D(instruction[10]), .Z(n16245)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_4_lut_adj_83.init = 16'h0008;
    LUT4 i17632_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22231), .B(n7762), .C(n22229), 
         .D(n22230), .Z(n17906)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17632_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hccc8;
    LUT4 i17682_2_lut_2_lut (.A(instruction[13]), .B(instruction[16]), .Z(n11804)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i17682_2_lut_2_lut.init = 16'h1111;
    LUT4 i5938_2_lut_4_lut (.A(instruction[10]), .B(instruction[11]), .C(instruction[9]), 
         .D(n8789), .Z(n7052)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i5938_2_lut_4_lut.init = 16'h0200;
    LUT4 i33_4_lut_3_lut (.A(instruction[12]), .B(instruction[14]), .C(instruction[15]), 
         .Z(n20)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+(C)))) */ ;
    defparam i33_4_lut_3_lut.init = 16'h2929;
    LUT4 i5926_2_lut_4_lut (.A(instruction[10]), .B(instruction[11]), .C(instruction[9]), 
         .D(n8789), .Z(n7080)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i5926_2_lut_4_lut.init = 16'h2000;
    LUT4 i2_2_lut_3_lut (.A(instruction[13]), .B(instruction[16]), .C(instruction[17]), 
         .Z(n7_adj_837)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i2_2_lut_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_4_lut_adj_84 (.A(instruction[9]), .B(n8789), .C(instruction[11]), 
         .D(instruction[10]), .Z(n16354)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_4_lut_adj_84.init = 16'h0040;
    LUT4 PrioSelect_585_i8_4_lut (.A(n6_adj_838), .B(n14_adj_711), .C(n7923), 
         .D(n7919), .Z(n8_adj_839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_585_i8_4_lut.init = 16'hcfca;
    LUT4 i1_2_lut_3_lut_adj_85 (.A(instruction[15]), .B(instruction[16]), 
         .C(instruction[17]), .Z(n16487)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(216[16:21])
    defparam i1_2_lut_3_lut_adj_85.init = 16'hfbfb;
    LUT4 i1_2_lut_4_lut_adj_86 (.A(instruction[9]), .B(n8789), .C(instruction[11]), 
         .D(instruction[10]), .Z(n16356)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_4_lut_adj_86.init = 16'h0080;
    LUT4 i16628_3_lut (.A(s_14_0), .B(s_15_0), .C(instruction[8]), .Z(n19798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16628_3_lut.init = 16'hcaca;
    LUT4 i16627_3_lut (.A(s_12_0), .B(s_13_0), .C(instruction[8]), .Z(n19797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16627_3_lut.init = 16'hcaca;
    LUT4 i16625_3_lut (.A(s_10_0), .B(s_11_0), .C(instruction[8]), .Z(n19795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16625_3_lut.init = 16'hcaca;
    PFUMX PrioSelect_137_i16 (.BLUT(n14_adj_840), .ALUT(n15_adj_841), .C0(n16998), 
          .Z(n16_adj_842)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i2_4_lut (.A(n16389), .B(n16_adj_843), .C(n13_adj_844), .D(C_N_342[8]), 
         .Z(n16391)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i2_4_lut.init = 16'ha080;
    LUT4 i16624_3_lut (.A(s_8_0), .B(s_9_0), .C(instruction[8]), .Z(n19794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16624_3_lut.init = 16'hcaca;
    LUT4 i16622_3_lut (.A(s_10_3), .B(s_11_3), .C(instruction[8]), .Z(n19792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16622_3_lut.init = 16'hcaca;
    LUT4 i16621_3_lut (.A(s_8_3), .B(s_9_3), .C(instruction[8]), .Z(n19791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16621_3_lut.init = 16'hcaca;
    LUT4 i16619_3_lut (.A(s_14_3), .B(s_15_3), .C(instruction[8]), .Z(n19789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16619_3_lut.init = 16'hcaca;
    LUT4 i16618_3_lut (.A(s_12_3), .B(s_13_3), .C(instruction[8]), .Z(n19788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16618_3_lut.init = 16'hcaca;
    LUT4 i44_4_lut_then_4_lut (.A(instruction[13]), .B(instruction[16]), 
         .C(instruction[14]), .D(C), .Z(n22318)) /* synthesis lut_function=(!(((C (D)+!C !(D))+!B)+!A)) */ ;
    defparam i44_4_lut_then_4_lut.init = 16'h0880;
    LUT4 i16616_3_lut (.A(s_10_4), .B(s_11_4), .C(instruction[8]), .Z(n19786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16616_3_lut.init = 16'hcaca;
    PFUMX PrioSelect_137_i13 (.BLUT(n8_adj_845), .ALUT(n12_adj_846), .C0(n16986), 
          .Z(n13_adj_847)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i16615_3_lut (.A(s_8_4), .B(s_9_4), .C(instruction[8]), .Z(n19785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16615_3_lut.init = 16'hcaca;
    LUT4 i16607_3_lut (.A(s_14_6), .B(s_15_6), .C(instruction[4]), .Z(n19777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16607_3_lut.init = 16'hcaca;
    LUT4 i16606_3_lut (.A(s_12_6), .B(s_13_6), .C(instruction[4]), .Z(n19776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16606_3_lut.init = 16'hcaca;
    LUT4 i16605_3_lut (.A(s_10_6), .B(s_11_6), .C(instruction[4]), .Z(n19775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16605_3_lut.init = 16'hcaca;
    LUT4 i16604_3_lut (.A(s_8_6), .B(s_9_6), .C(instruction[4]), .Z(n19774)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16604_3_lut.init = 16'hcaca;
    LUT4 i16603_3_lut (.A(s_6_6), .B(s_7_6), .C(instruction[4]), .Z(n19773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16603_3_lut.init = 16'hcaca;
    LUT4 i44_4_lut_else_4_lut (.A(Z), .B(instruction[13]), .C(instruction[16]), 
         .D(instruction[14]), .Z(n22317)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam i44_4_lut_else_4_lut.init = 16'h400f;
    LUT4 i8_4_lut (.A(Z_N_367[6]), .B(n16_adj_848), .C(n16524), .D(Z_N_367[2]), 
         .Z(n14780)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i8_4_lut.init = 16'h0004;
    LUT4 i16602_3_lut (.A(s_4_6), .B(s_5_6), .C(instruction[4]), .Z(n19772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16602_3_lut.init = 16'hcaca;
    LUT4 i16601_3_lut (.A(s_2_6), .B(s_3_6), .C(instruction[4]), .Z(n19771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16601_3_lut.init = 16'hcaca;
    LUT4 i16600_3_lut (.A(s_0_6), .B(s_1_6), .C(instruction[4]), .Z(n19770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16600_3_lut.init = 16'hcaca;
    LUT4 i16598_3_lut (.A(s_14_4), .B(s_15_4), .C(instruction[8]), .Z(n19768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16598_3_lut.init = 16'hcaca;
    LUT4 i8920_2_lut_3_lut (.A(instruction[12]), .B(instruction[14]), .C(instruction[13]), 
         .Z(n8_adj_849)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i8920_2_lut_3_lut.init = 16'hfefe;
    LUT4 i16597_3_lut (.A(s_12_4), .B(s_13_4), .C(instruction[8]), .Z(n19767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16597_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_77_i4_4_lut (.A(n2), .B(C), .C(n16261), .D(n16252), 
         .Z(n4_adj_850)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_77_i4_4_lut.init = 16'hc0ca;
    LUT4 i16595_3_lut (.A(s_10_5), .B(s_11_5), .C(instruction[8]), .Z(n19765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16595_3_lut.init = 16'hcaca;
    PFUMX PrioSelect_133_i19 (.BLUT(n15_adj_752), .ALUT(n17_adj_851), .C0(n16969), 
          .Z(n455)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i16594_3_lut (.A(s_8_5), .B(s_9_5), .C(instruction[8]), .Z(n19764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16594_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_87 (.A(instruction[9]), .B(n8789), .C(instruction[10]), 
         .D(instruction[11]), .Z(n6886)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_4_lut_adj_87.init = 16'h4000;
    LUT4 PrioSelect_105_i8_4_lut (.A(n6_adj_852), .B(n7_adj_473), .C(n16268), 
         .D(n16284), .Z(n8_adj_853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_105_i8_4_lut.init = 16'hcfca;
    LUT4 i16592_3_lut (.A(s_14_5), .B(s_15_5), .C(instruction[8]), .Z(n19762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16592_3_lut.init = 16'hcaca;
    LUT4 i16591_3_lut (.A(s_12_5), .B(s_13_5), .C(instruction[8]), .Z(n19761)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16591_3_lut.init = 16'hcaca;
    PFUMX PrioSelect_129_i19 (.BLUT(n15_adj_772), .ALUT(n17_adj_854), .C0(n16969), 
          .Z(n451)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i16589_3_lut (.A(s_10_6), .B(s_11_6), .C(instruction[8]), .Z(n19759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16589_3_lut.init = 16'hcaca;
    LUT4 i16588_3_lut (.A(s_8_6), .B(s_9_6), .C(instruction[8]), .Z(n19758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16588_3_lut.init = 16'hcaca;
    LUT4 i16586_3_lut (.A(s_14_6), .B(s_15_6), .C(instruction[8]), .Z(n19756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16586_3_lut.init = 16'hcaca;
    LUT4 i16585_3_lut (.A(s_12_6), .B(s_13_6), .C(instruction[8]), .Z(n19755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16585_3_lut.init = 16'hcaca;
    LUT4 i17551_2_lut (.A(n9164), .B(n20152), .Z(n16685)) /* synthesis lut_function=(A+(B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17551_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_515_3_lut (.A(n2075), .B(instruction[8]), .C(instruction[9]), 
         .Z(n22082)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(223[39:43])
    defparam i1_2_lut_rep_515_3_lut.init = 16'h0202;
    LUT4 i16583_3_lut (.A(s_10_7), .B(s_11_7), .C(instruction[8]), .Z(n19753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16583_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_88 (.A(instruction[15]), .B(instruction[16]), 
         .C(instruction[17]), .Z(n10_adj_698)) /* synthesis lut_function=((B+(C))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[16:28])
    defparam i1_2_lut_3_lut_adj_88.init = 16'hfdfd;
    LUT4 i16582_3_lut (.A(s_8_7), .B(s_9_7), .C(instruction[8]), .Z(n19752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16582_3_lut.init = 16'hcaca;
    LUT4 i16580_3_lut (.A(s_14_7), .B(s_15_7), .C(instruction[8]), .Z(n19750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16580_3_lut.init = 16'hcaca;
    LUT4 i16579_3_lut (.A(s_12_7), .B(s_13_7), .C(instruction[8]), .Z(n19749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16579_3_lut.init = 16'hcaca;
    LUT4 i16577_3_lut (.A(s_10_1), .B(s_11_1), .C(instruction[8]), .Z(n19747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16577_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_109_i4_4_lut (.A(n2_adj_855), .B(C), .C(n16277), .D(n16259), 
         .Z(n4_adj_856)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_109_i4_4_lut.init = 16'hc0ca;
    LUT4 i16576_3_lut (.A(s_8_1), .B(s_9_1), .C(instruction[8]), .Z(n19746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16576_3_lut.init = 16'hcaca;
    LUT4 i16574_3_lut (.A(s_14_1), .B(s_15_1), .C(instruction[8]), .Z(n19744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16574_3_lut.init = 16'hcaca;
    LUT4 i17627_2_lut_2_lut (.A(instruction[16]), .B(instruction[15]), .Z(n16618)) /* synthesis lut_function=((B)+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i17627_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_89 (.A(n22304), .B(n22284), .C(n7746), 
         .D(n22307), .Z(n1[19])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_89.init = 16'h0080;
    LUT4 i17215_3_lut_4_lut (.A(n22153), .B(n22087), .C(n14_adj_857), 
         .D(n10_adj_858), .Z(n15_adj_665)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17215_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16573_3_lut (.A(s_12_1), .B(s_13_1), .C(instruction[8]), .Z(n19743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16573_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_90 (.A(instruction[10]), .B(instruction[11]), 
         .C(instruction[8]), .D(instruction[9]), .Z(n16375)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam i1_2_lut_4_lut_adj_90.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_91 (.A(n22304), .B(n22284), .C(n22282), 
         .D(n22307), .Z(n1[15])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_91.init = 16'h8000;
    LUT4 PrioSelect_297_i12_3_lut_4_lut (.A(n22231), .B(n7762), .C(Z_N_378[7]), 
         .D(n11_adj_828), .Z(n12_adj_859)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_297_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_269_i12_3_lut_4_lut (.A(n22231), .B(n7762), .C(Z_N_378[0]), 
         .D(n11_adj_834), .Z(n12_adj_860)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_269_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_3_lut_4_lut_adj_92 (.A(instruction[12]), .B(instruction[15]), 
         .C(instruction[14]), .D(n5_adj_861), .Z(n14428)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;
    defparam i2_3_lut_4_lut_adj_92.init = 16'h5400;
    LUT4 i1_2_lut_3_lut_adj_93 (.A(instruction[15]), .B(instruction[16]), 
         .C(instruction[17]), .Z(n10_adj_586)) /* synthesis lut_function=(A+(B+(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[16:28])
    defparam i1_2_lut_3_lut_adj_93.init = 16'hfefe;
    LUT4 i1_2_lut_adj_94 (.A(instruction[13]), .B(instruction[16]), .Z(n5_adj_861)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_2_lut_adj_94.init = 16'h8888;
    PFUMX PrioSelect_125_i19 (.BLUT(n15_adj_762), .ALUT(n17_adj_862), .C0(n16969), 
          .Z(n447)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_3_lut_adj_95 (.A(instruction[12]), .B(instruction[14]), 
         .C(instruction[13]), .Z(n8_adj_695)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(240[16:24])
    defparam i1_2_lut_3_lut_adj_95.init = 16'hdfdf;
    LUT4 i6099_2_lut_3_lut_4_lut (.A(n160), .B(n7646), .C(instruction[3]), 
         .D(instruction[8]), .Z(n8789)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i6099_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 instruction_17__I_0_569_i10_2_lut_3_lut (.A(instruction[15]), .B(instruction[16]), 
         .C(instruction[17]), .Z(n10_adj_863)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[17:26])
    defparam instruction_17__I_0_569_i10_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut_adj_96 (.A(instruction[12]), .B(instruction[14]), 
         .C(instruction[13]), .Z(n8_adj_708)) /* synthesis lut_function=((B+(C))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(234[16:28])
    defparam i1_2_lut_3_lut_adj_96.init = 16'hfdfd;
    LUT4 n8_bdd_2_lut_3_lut_4_lut (.A(instruction[12]), .B(instruction[14]), 
         .C(instruction[13]), .D(instruction[16]), .Z(n21531)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam n8_bdd_2_lut_3_lut_4_lut.init = 16'hffdf;
    LUT4 i1_4_lut_4_lut (.A(instruction[12]), .B(Z), .C(n21796), .D(n7628), 
         .Z(n19)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_4_lut_4_lut.init = 16'h5044;
    LUT4 PrioSelect_233_i9_3_lut_4_lut (.A(n22101), .B(n7762), .C(n7_adj_500), 
         .D(C), .Z(n9_adj_864)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_233_i9_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_121_i19 (.BLUT(n15_adj_769), .ALUT(n17_adj_865), .C0(n16969), 
          .Z(n443)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i2_3_lut_4_lut_adj_97 (.A(n14802), .B(instruction[15]), .C(instruction[14]), 
         .D(instruction[12]), .Z(n14803)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_4_lut_adj_97.init = 16'h0020;
    LUT4 i17236_3_lut_4_lut (.A(n22159), .B(n22088), .C(n14_adj_726), 
         .D(n10_adj_866), .Z(n15_adj_621)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17236_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17226_3_lut_4_lut (.A(n22159), .B(n22088), .C(n14_adj_697), 
         .D(n10_adj_867), .Z(n15_adj_637)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17226_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17232_3_lut_4_lut (.A(n22159), .B(n22088), .C(n14_adj_715), 
         .D(n10_adj_868), .Z(n15_adj_629)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17232_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17230_3_lut_4_lut (.A(n22159), .B(n22088), .C(n14_adj_704), 
         .D(n10_adj_869), .Z(n15_adj_633)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17230_3_lut_4_lut.init = 16'hf1e0;
    PFUMX PrioSelect_117_i19 (.BLUT(n15_adj_775), .ALUT(n17_adj_870), .C0(n16969), 
          .Z(n439)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17479_4_lut (.A(Z_N_378[0]), .B(n20080), .C(n10_adj_871), .D(Z_N_378[6]), 
         .Z(Z_N_377)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[119:138])
    defparam i17479_4_lut.init = 16'h0004;
    LUT4 i17478_4_lut (.A(Z_N_378[3]), .B(Z_N_378[1]), .C(Z_N_378[5]), 
         .D(Z_N_378[7]), .Z(n20080)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[119:138])
    defparam i17478_4_lut.init = 16'h0001;
    LUT4 i2_2_lut (.A(Z_N_378[2]), .B(Z_N_378[4]), .Z(n10_adj_871)) /* synthesis lut_function=(A+(B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[119:138])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 instruction_17__I_0_562_i11_2_lut_3_lut_4_lut (.A(instruction[12]), 
         .B(instruction[14]), .C(instruction[13]), .D(n10_adj_776), .Z(n11_adj_872)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(299[17:21])
    defparam instruction_17__I_0_562_i11_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i17234_3_lut_4_lut (.A(n22159), .B(n22088), .C(n14_adj_718), 
         .D(n10_adj_873), .Z(n15_adj_627)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17234_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17228_3_lut_4_lut (.A(n22159), .B(n22088), .C(n14_adj_700), 
         .D(n10_adj_874), .Z(n15_adj_635)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17228_3_lut_4_lut.init = 16'hf1e0;
    PFUMX PrioSelect_113_i19 (.BLUT(n15_adj_759), .ALUT(n17_adj_875), .C0(n16969), 
          .Z(n435)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_265_i9_3_lut_4_lut (.A(n22093), .B(n7762), .C(n7_adj_500), 
         .D(C), .Z(n9_adj_876)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_265_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i17250_3_lut_4_lut (.A(n22165), .B(n22089), .C(n14_adj_877), 
         .D(n10_adj_878), .Z(n15_adj_600)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17250_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16571_3_lut (.A(s_10_2), .B(s_11_2), .C(instruction[8]), .Z(n19741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16571_3_lut.init = 16'hcaca;
    LUT4 i16570_3_lut (.A(s_8_2), .B(s_9_2), .C(instruction[8]), .Z(n19740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16570_3_lut.init = 16'hcaca;
    PFUMX PrioSelect_105_i16 (.BLUT(n14_adj_653), .ALUT(n15), .C0(n16814), 
          .Z(n16_adj_879)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_141_i4_4_lut (.A(n2_adj_880), .B(C), .C(n16260), .D(n16244), 
         .Z(n4_adj_881)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_141_i4_4_lut.init = 16'hc0ca;
    LUT4 i16568_3_lut (.A(s_14_2), .B(s_15_2), .C(instruction[8]), .Z(n19738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16568_3_lut.init = 16'hcaca;
    LUT4 i16567_3_lut (.A(s_12_2), .B(s_13_2), .C(instruction[8]), .Z(n19737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16567_3_lut.init = 16'hcaca;
    LUT4 i16563_3_lut (.A(s_6_0), .B(s_7_0), .C(instruction[8]), .Z(n19733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16563_3_lut.init = 16'hcaca;
    LUT4 i17240_3_lut_4_lut (.A(n22165), .B(n22089), .C(n14_adj_882), 
         .D(n10_adj_883), .Z(n15_adj_612)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17240_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16562_3_lut (.A(s_4_0), .B(s_5_0), .C(instruction[8]), .Z(n19732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16562_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_169_i8_4_lut (.A(n6_adj_884), .B(n7_adj_473), .C(n16269), 
         .D(n16285), .Z(n8_adj_885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_169_i8_4_lut.init = 16'hcfca;
    LUT4 i16561_3_lut (.A(s_2_0), .B(s_3_0), .C(instruction[8]), .Z(n19731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16561_3_lut.init = 16'hcaca;
    LUT4 i17246_3_lut_4_lut (.A(n22165), .B(n22089), .C(n14_adj_886), 
         .D(n10_adj_887), .Z(n15_adj_605)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17246_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16560_3_lut (.A(s_0_0), .B(s_1_0), .C(instruction[8]), .Z(n19730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16560_3_lut.init = 16'hcaca;
    LUT4 i16556_3_lut (.A(s_6_3), .B(s_7_3), .C(instruction[8]), .Z(n19726)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16556_3_lut.init = 16'hcaca;
    LUT4 i16555_3_lut (.A(s_4_3), .B(s_5_3), .C(instruction[8]), .Z(n19725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16555_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_269_i15_3_lut_4_lut (.A(n22232), .B(n7762), .C(n1108[0]), 
         .D(n5_adj_602), .Z(n15_adj_888)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_269_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i16554_3_lut (.A(s_2_3), .B(s_3_3), .C(instruction[8]), .Z(n19724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16554_3_lut.init = 16'hcaca;
    LUT4 i16553_3_lut (.A(s_0_3), .B(s_1_3), .C(instruction[8]), .Z(n19723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16553_3_lut.init = 16'hcaca;
    PFUMX PrioSelect_101_i19 (.BLUT(n15_adj_889), .ALUT(n17_adj_890), .C0(n16685), 
          .Z(n423)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i16549_3_lut (.A(s_6_4), .B(s_7_4), .C(instruction[8]), .Z(n19719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16549_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_173_i4_4_lut (.A(n2_adj_891), .B(C), .C(n16276), .D(n16258), 
         .Z(n4_adj_892)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_173_i4_4_lut.init = 16'hc0ca;
    LUT4 i16548_3_lut (.A(s_4_4), .B(s_5_4), .C(instruction[8]), .Z(n19718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16548_3_lut.init = 16'hcaca;
    LUT4 i16547_3_lut (.A(s_2_4), .B(s_3_4), .C(instruction[8]), .Z(n19717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16547_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_293_i12_3_lut_4_lut (.A(n22232), .B(n7762), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_893)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_293_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17244_3_lut_4_lut (.A(n22165), .B(n22089), .C(n14_adj_894), 
         .D(n10_adj_895), .Z(n15_adj_607)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17244_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_289_i12_3_lut_4_lut (.A(n22232), .B(n7762), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_896)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_289_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i16546_3_lut (.A(s_0_4), .B(s_1_4), .C(instruction[8]), .Z(n19716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16546_3_lut.init = 16'hcaca;
    LUT4 i17248_3_lut_4_lut (.A(n22165), .B(n22089), .C(n14_adj_897), 
         .D(n10_adj_898), .Z(n15_adj_603)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17248_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17242_3_lut_4_lut (.A(n22165), .B(n22089), .C(n14_adj_899), 
         .D(n10_adj_900), .Z(n15_adj_610)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17242_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16542_3_lut (.A(s_6_5), .B(s_7_5), .C(instruction[8]), .Z(n19712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16542_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_205_i4_4_lut (.A(n2_adj_901), .B(C), .C(n83), .D(n54[4]), 
         .Z(n4_adj_902)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_205_i4_4_lut.init = 16'hc0ca;
    PFUMX PrioSelect_97_i19 (.BLUT(n15_adj_903), .ALUT(n17_adj_904), .C0(n16685), 
          .Z(n419)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_297_i9_3_lut_4_lut (.A(n22095), .B(n7762), .C(n7_adj_500), 
         .D(C), .Z(n9_adj_905)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_297_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i16541_3_lut (.A(s_4_5), .B(s_5_5), .C(instruction[8]), .Z(n19711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16541_3_lut.init = 16'hcaca;
    LUT4 i17263_3_lut_4_lut (.A(n22171), .B(n22090), .C(n14_adj_906), 
         .D(n10_adj_907), .Z(n15_adj_581)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17263_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_285_i12_3_lut_4_lut (.A(n22232), .B(n7762), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_908)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_285_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_281_i12_3_lut_4_lut (.A(n22232), .B(n7762), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_909)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_281_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17253_3_lut_4_lut (.A(n22171), .B(n22090), .C(n14_adj_910), 
         .D(n10_adj_911), .Z(n15_adj_594)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17253_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17259_3_lut_4_lut (.A(n22171), .B(n22090), .C(n14_adj_912), 
         .D(n10_adj_913), .Z(n15_adj_587)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17259_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_233_i8_4_lut (.A(n6_adj_914), .B(n7_adj_473), .C(n151[4]), 
         .D(n146), .Z(n8_adj_915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_233_i8_4_lut.init = 16'hcfca;
    LUT4 i16540_3_lut (.A(s_2_5), .B(s_3_5), .C(instruction[8]), .Z(n19710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16540_3_lut.init = 16'hcaca;
    LUT4 i16539_3_lut (.A(s_0_5), .B(s_1_5), .C(instruction[8]), .Z(n19709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16539_3_lut.init = 16'hcaca;
    PFUMX PrioSelect_93_i19 (.BLUT(n15_adj_916), .ALUT(n17_adj_917), .C0(n16685), 
          .Z(n415)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i16535_3_lut (.A(s_6_7), .B(s_7_7), .C(instruction[8]), .Z(n19705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16535_3_lut.init = 16'hcaca;
    LUT4 i5932_2_lut_3_lut_4_lut (.A(n160), .B(n16421), .C(n7762), .D(n7726), 
         .Z(n7066)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i5932_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_98 (.A(n160), .B(n16421), .C(n11714), 
         .D(n7876), .Z(n16246)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_3_lut_4_lut_adj_98.init = 16'h0800;
    LUT4 PrioSelect_277_i12_3_lut_4_lut (.A(n22232), .B(n7762), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_918)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_277_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_273_i12_3_lut_4_lut (.A(n22232), .B(n7762), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_919)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_273_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_99 (.A(n160), .B(n16421), .C(n11714), 
         .D(n7726), .Z(n16251)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_3_lut_4_lut_adj_99.init = 16'h0800;
    LUT4 i17257_3_lut_4_lut (.A(n22171), .B(n22090), .C(n14_adj_920), 
         .D(n10_adj_921), .Z(n15_adj_589)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17257_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_297_i15_3_lut_4_lut (.A(n22232), .B(n7762), .C(n1108[7]), 
         .D(n9_adj_905), .Z(n15_adj_598)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_297_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_237_i4_4_lut (.A(n2_adj_922), .B(C), .C(n82), .D(n54[5]), 
         .Z(n4_adj_923)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_237_i4_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_adj_100 (.A(instruction[8]), .B(instruction[9]), .Z(n7726)) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(225[39:43])
    defparam i1_2_lut_adj_100.init = 16'h2222;
    PFUMX PrioSelect_89_i19 (.BLUT(n15_adj_924), .ALUT(n17_adj_925), .C0(n16685), 
          .Z(n411)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 n2083_bdd_4_lut_17862 (.A(n22109), .B(n2085), .C(n16312), .D(n16392), 
         .Z(n21115)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam n2083_bdd_4_lut_17862.init = 16'h1fff;
    LUT4 i16534_3_lut (.A(s_4_7), .B(s_5_7), .C(instruction[8]), .Z(n19704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16534_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_297_i10_3_lut_4_lut (.A(n22233), .B(n7762), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_926)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_297_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_269_i4_4_lut (.A(n2_adj_927), .B(C), .C(n81), .D(n54[6]), 
         .Z(n4_adj_928)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_269_i4_4_lut.init = 16'hc0ca;
    LUT4 i17261_3_lut_4_lut (.A(n22171), .B(n22090), .C(n14_adj_929), 
         .D(n10_adj_930), .Z(n15_adj_584)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17261_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16533_3_lut (.A(s_2_7), .B(s_3_7), .C(instruction[8]), .Z(n19703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16533_3_lut.init = 16'hcaca;
    LUT4 i16532_3_lut (.A(s_0_7), .B(s_1_7), .C(instruction[8]), .Z(n19702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16532_3_lut.init = 16'hcaca;
    LUT4 i16528_3_lut (.A(s_6_6), .B(s_7_6), .C(instruction[8]), .Z(n19698)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16528_3_lut.init = 16'hcaca;
    LUT4 i16527_3_lut (.A(s_4_6), .B(s_5_6), .C(instruction[8]), .Z(n19697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16527_3_lut.init = 16'hcaca;
    LUT4 i17255_3_lut_4_lut (.A(n22171), .B(n22090), .C(n14_adj_931), 
         .D(n10_adj_932), .Z(n15_adj_591)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17255_3_lut_4_lut.init = 16'hf1e0;
    PFUMX PrioSelect_85_i19 (.BLUT(n15_adj_933), .ALUT(n17_adj_934), .C0(n16685), 
          .Z(n407)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i3_4_lut_then_4_lut (.A(instruction[17]), .B(instruction[12]), 
         .C(instruction[13]), .D(instruction[14]), .Z(n22321)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i3_4_lut_then_4_lut.init = 16'hdfff;
    LUT4 PrioSelect_297_i8_4_lut (.A(n6_adj_935), .B(n7_adj_473), .C(n151[6]), 
         .D(n143), .Z(n8_adj_936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_297_i8_4_lut.init = 16'hcfca;
    LUT4 i2138_3_lut_4_lut (.A(n22233), .B(n7762), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_937)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i2138_3_lut_4_lut.init = 16'hf780;
    LUT4 i16526_3_lut (.A(s_2_6), .B(s_3_6), .C(instruction[8]), .Z(n19696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16526_3_lut.init = 16'hcaca;
    LUT4 i16525_3_lut (.A(s_0_6), .B(s_1_6), .C(instruction[8]), .Z(n19695)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16525_3_lut.init = 16'hcaca;
    LUT4 i16521_3_lut (.A(s_6_1), .B(s_7_1), .C(instruction[8]), .Z(n19691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16521_3_lut.init = 16'hcaca;
    LUT4 i16520_3_lut (.A(s_4_1), .B(s_5_1), .C(instruction[8]), .Z(n19690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16520_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut_else_4_lut (.A(instruction[15]), .B(instruction[17]), 
         .C(instruction[12]), .D(instruction[13]), .Z(n22320)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i3_4_lut_else_4_lut.init = 16'hfff7;
    LUT4 i16519_3_lut (.A(s_2_1), .B(s_3_1), .C(instruction[8]), .Z(n19689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16519_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_301_i4_4_lut (.A(n2_adj_938), .B(C), .C(n80), .D(n54[7]), 
         .Z(n4_adj_939)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_301_i4_4_lut.init = 16'hc0ca;
    LUT4 i16518_3_lut (.A(s_0_1), .B(s_1_1), .C(instruction[8]), .Z(n19688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16518_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_293_i13_3_lut_4_lut (.A(n22233), .B(n7762), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_940)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_293_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 instruction_17__I_0_554_i9_2_lut (.A(instruction[16]), .B(instruction[17]), 
         .Z(n9_adj_707)) /* synthesis lut_function=((B)+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(216[16:21])
    defparam instruction_17__I_0_554_i9_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_adj_101 (.A(instruction[14]), .B(instruction[13]), .Z(n8050)) /* synthesis lut_function=(A+(B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_2_lut_adj_101.init = 16'heeee;
    LUT4 i16514_3_lut (.A(s_6_2), .B(s_7_2), .C(instruction[8]), .Z(n19684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16514_3_lut.init = 16'hcaca;
    LUT4 i16513_3_lut (.A(s_4_2), .B(s_5_2), .C(instruction[8]), .Z(n19683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16513_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_333_i4_4_lut (.A(n2_adj_941), .B(C), .C(n16351), .D(n16347), 
         .Z(n4_adj_942)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_333_i4_4_lut.init = 16'hc0ca;
    PFUMX PrioSelect_81_i19 (.BLUT(n15_adj_943), .ALUT(n17_adj_944), .C0(n16685), 
          .Z(n403)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i16512_3_lut (.A(s_2_2), .B(s_3_2), .C(instruction[8]), .Z(n19682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16512_3_lut.init = 16'hcaca;
    LUT4 i16511_3_lut (.A(s_0_2), .B(s_1_2), .C(instruction[8]), .Z(n19681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16511_3_lut.init = 16'hcaca;
    LUT4 i16503_3_lut (.A(s_14_0), .B(s_15_0), .C(instruction[4]), .Z(n19673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16503_3_lut.init = 16'hcaca;
    LUT4 i16502_3_lut (.A(s_12_0), .B(s_13_0), .C(instruction[4]), .Z(n19672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16502_3_lut.init = 16'hcaca;
    LUT4 i16501_3_lut (.A(s_10_0), .B(s_11_0), .C(instruction[4]), .Z(n19671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16501_3_lut.init = 16'hcaca;
    LUT4 i16500_3_lut (.A(s_8_0), .B(s_9_0), .C(instruction[4]), .Z(n19670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16500_3_lut.init = 16'hcaca;
    LUT4 i16499_3_lut (.A(s_6_0), .B(s_7_0), .C(instruction[4]), .Z(n19669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16499_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_102 (.A(n160), .B(n16421), .C(n7908), 
         .D(n7726), .Z(n6900)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_3_lut_4_lut_adj_102.init = 16'h8000;
    LUT4 PrioSelect_361_i8_4_lut (.A(n6_adj_945), .B(n14_adj_711), .C(n16341), 
         .D(n16327), .Z(n8_adj_946)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_361_i8_4_lut.init = 16'hcfca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_103 (.A(n160), .B(n16421), .C(n16312), 
         .D(n7876), .Z(n16358)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_3_lut_4_lut_adj_103.init = 16'h8000;
    PFUMX i119 (.BLUT(n14358), .ALUT(n7696), .C0(instruction[17]), .Z(n61));
    LUT4 i1_2_lut_3_lut_4_lut_adj_104 (.A(n22304), .B(n22284), .C(n22285), 
         .D(n22307), .Z(n1[7])) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_104.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_105 (.A(n160), .B(n16421), .C(n16312), 
         .D(n7726), .Z(n16357)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_3_lut_4_lut_adj_105.init = 16'h8000;
    LUT4 i16498_3_lut (.A(s_4_0), .B(s_5_0), .C(instruction[4]), .Z(n19668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16498_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_365_i4_4_lut (.A(n2_adj_947), .B(C), .C(n16316), .D(n16350), 
         .Z(n4_adj_948)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_365_i4_4_lut.init = 16'hc0ca;
    LUT4 i16497_3_lut (.A(s_2_0), .B(s_3_0), .C(instruction[4]), .Z(n19667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16497_3_lut.init = 16'hcaca;
    LUT4 i16496_3_lut (.A(s_0_0), .B(s_1_0), .C(instruction[4]), .Z(n19666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16496_3_lut.init = 16'hcaca;
    LUT4 i16488_3_lut (.A(s_14_1), .B(s_15_1), .C(instruction[4]), .Z(n19658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16488_3_lut.init = 16'hcaca;
    LUT4 i16487_3_lut (.A(s_12_1), .B(s_13_1), .C(instruction[4]), .Z(n19657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16487_3_lut.init = 16'hcaca;
    LUT4 i16486_3_lut (.A(s_10_1), .B(s_11_1), .C(instruction[4]), .Z(n19656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16486_3_lut.init = 16'hcaca;
    LUT4 i16485_3_lut (.A(s_8_1), .B(s_9_1), .C(instruction[4]), .Z(n19655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16485_3_lut.init = 16'hcaca;
    LUT4 i16484_3_lut (.A(s_6_1), .B(s_7_1), .C(instruction[4]), .Z(n19654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16484_3_lut.init = 16'hcaca;
    LUT4 i16483_3_lut (.A(s_4_1), .B(s_5_1), .C(instruction[4]), .Z(n19653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16483_3_lut.init = 16'hcaca;
    LUT4 i16482_3_lut (.A(s_2_1), .B(s_3_1), .C(instruction[4]), .Z(n19652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16482_3_lut.init = 16'hcaca;
    LUT4 i16481_3_lut (.A(s_0_1), .B(s_1_1), .C(instruction[4]), .Z(n19651)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16481_3_lut.init = 16'hcaca;
    LUT4 i16473_3_lut (.A(s_14_5), .B(s_15_5), .C(instruction[4]), .Z(n19643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16473_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_397_i4_4_lut (.A(n2_adj_949), .B(C), .C(n16348), .D(n16355), 
         .Z(n4_adj_950)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_397_i4_4_lut.init = 16'hc0ca;
    LUT4 i16472_3_lut (.A(s_12_5), .B(s_13_5), .C(instruction[4]), .Z(n19642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16472_3_lut.init = 16'hcaca;
    PFUMX PrioSelect_461_i16 (.BLUT(n14_adj_951), .ALUT(n15_adj_952), .C0(n19022), 
          .Z(n16_adj_953)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i16471_3_lut (.A(s_10_5), .B(s_11_5), .C(instruction[4]), .Z(n19641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16471_3_lut.init = 16'hcaca;
    LUT4 i16470_3_lut (.A(s_8_5), .B(s_9_5), .C(instruction[4]), .Z(n19640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16470_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_289_i13_3_lut_4_lut (.A(n22233), .B(n7762), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_954)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_289_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_285_i13_3_lut_4_lut (.A(n22233), .B(n7762), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_955)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_285_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 n8932_bdd_4_lut (.A(n1339), .B(n1341), .C(clk_in_c_enable_115), 
         .D(clk_in_c_enable_109), .Z(n21515)) /* synthesis lut_function=(A+!(B ((D)+!C))) */ ;
    defparam n8932_bdd_4_lut.init = 16'hbbfb;
    LUT4 PrioSelect_329_i9_3_lut_4_lut (.A(n22097), .B(n7762), .C(n7_adj_500), 
         .D(C), .Z(n9_adj_956)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_329_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_281_i13_3_lut_4_lut (.A(n22233), .B(n7762), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_957)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_281_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i5920_2_lut_3_lut_4_lut (.A(n160), .B(n16421), .C(n7762), .D(n7876), 
         .Z(n7094)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i5920_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 PrioSelect_425_i8_4_lut (.A(n6_adj_958), .B(n14_adj_711), .C(n16338), 
         .D(n16332), .Z(n8_adj_959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_425_i8_4_lut.init = 16'hcfca;
    PFUMX PrioSelect_397_i16 (.BLUT(n14_adj_960), .ALUT(n15_adj_961), .C0(n18654), 
          .Z(n16_adj_962)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_277_i13_3_lut_4_lut (.A(n22233), .B(n7762), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_963)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_277_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i17675_2_lut_rep_514 (.A(rst_n_in), .B(n5_adj_964), .Z(clk_in_c_enable_175)) /* synthesis lut_function=(!(A (B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i17675_2_lut_rep_514.init = 16'h7777;
    PFUMX PrioSelect_333_i16 (.BLUT(n14_adj_965), .ALUT(n15_adj_966), .C0(n18286), 
          .Z(n16_adj_967)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 n8_bdd_4_lut_18613 (.A(n16484), .B(instruction[12]), .C(instruction[15]), 
         .D(instruction[16]), .Z(n21530)) /* synthesis lut_function=(A+(B+!(C (D)+!C !(D)))) */ ;
    defparam n8_bdd_4_lut_18613.init = 16'heffe;
    LUT4 seg_led_2_c_bdd_2_lut_18089_3_lut (.A(rst_n_in), .B(n5_adj_964), 
         .C(n21515), .Z(n21516)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam seg_led_2_c_bdd_2_lut_18089_3_lut.init = 16'h7070;
    PFUMX PrioSelect_269_i16 (.BLUT(n14_adj_968), .ALUT(n15_adj_888), .C0(n17918), 
          .Z(n16_adj_969)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_273_i13_3_lut_4_lut (.A(n22233), .B(n7762), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_970)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_273_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_429_i4_4_lut (.A(n2_adj_971), .B(C), .C(n16315), .D(n16349), 
         .Z(n4_adj_972)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_429_i4_4_lut.init = 16'hc0ca;
    PFUMX PrioSelect_205_i16 (.BLUT(n14_adj_973), .ALUT(n15_adj_974), .C0(n17550), 
          .Z(n16_adj_975)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17277_3_lut_4_lut (.A(n22177), .B(n22091), .C(n14_adj_976), 
         .D(n10_adj_712), .Z(n15_adj_561)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17277_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_106 (.A(n22304), .B(n22284), .C(n22285), 
         .D(n22307), .Z(n1[3])) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_106.init = 16'h0008;
    LUT4 i17267_3_lut_4_lut (.A(n22177), .B(n22091), .C(n14_adj_977), 
         .D(n10_adj_699), .Z(n15_adj_572)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17267_3_lut_4_lut.init = 16'hf1e0;
    PFUMX PrioSelect_141_i16 (.BLUT(n14_adj_978), .ALUT(n15_adj_979), .C0(n17182), 
          .Z(n16_adj_980)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17273_3_lut_4_lut (.A(n22177), .B(n22091), .C(n14_adj_981), 
         .D(n10_adj_706), .Z(n15_adj_566)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17273_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17583_2_lut_3_lut_4_lut (.A(n22264), .B(n7876), .C(n20184), 
         .D(n7908), .Z(n19421)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17583_2_lut_3_lut_4_lut.init = 16'hf4f0;
    PFUMX PrioSelect_77_i16 (.BLUT(n14_adj_649), .ALUT(n15_adj_982), .C0(n16814), 
          .Z(n16_adj_983)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_273_i14_3_lut_4_lut (.A(n22234), .B(n7762), .C(Z_N_387[1]), 
         .D(n13_adj_970), .Z(n14_adj_882)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_273_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_277_i14_3_lut_4_lut (.A(n22234), .B(n7762), .C(Z_N_387[2]), 
         .D(n13_adj_963), .Z(n14_adj_899)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_277_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX i118 (.BLUT(n29), .ALUT(n34), .C0(n24), .Z(n85));
    LUT4 PrioSelect_281_i14_3_lut_4_lut (.A(n22234), .B(n7762), .C(Z_N_387[3]), 
         .D(n13_adj_957), .Z(n14_adj_894)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_281_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_107 (.A(instruction[14]), .B(instruction[13]), .Z(n16484)) /* synthesis lut_function=(A+!(B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(240[16:24])
    defparam i1_2_lut_adj_107.init = 16'hbbbb;
    LUT4 i8208_4_lut (.A(n19928), .B(st_zc[3]), .C(n21), .D(st_zc[2]), 
         .Z(n30)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(376[66:84])
    defparam i8208_4_lut.init = 16'h3022;
    LUT4 i16469_3_lut (.A(s_6_5), .B(s_7_5), .C(instruction[4]), .Z(n19639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16469_3_lut.init = 16'hcaca;
    PFUMX PrioSelect_525_i16 (.BLUT(n14_adj_984), .ALUT(n15_adj_985), .C0(n19390), 
          .Z(n16_adj_986)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_285_i14_3_lut_4_lut (.A(n22234), .B(n7762), .C(Z_N_387[4]), 
         .D(n13_adj_955), .Z(n14_adj_886)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_285_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_289_i14_3_lut_4_lut (.A(n22234), .B(n7762), .C(Z_N_387[5]), 
         .D(n13_adj_954), .Z(n14_adj_897)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_289_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_493_i16 (.BLUT(n14_adj_987), .ALUT(n15_adj_624), .C0(n19206), 
          .Z(n16_adj_988)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_201_i12_3_lut_4_lut (.A(n22237), .B(n11714), .C(Z_N_378[7]), 
         .D(n11_adj_688), .Z(n12_adj_674)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_201_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i16468_3_lut (.A(s_4_5), .B(s_5_5), .C(instruction[4]), .Z(n19638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16468_3_lut.init = 16'hcaca;
    LUT4 i17271_3_lut_4_lut (.A(n22177), .B(n22091), .C(n14_adj_989), 
         .D(n10_adj_702), .Z(n15_adj_568)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17271_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17275_3_lut_4_lut (.A(n22177), .B(n22091), .C(n14_adj_990), 
         .D(n10_adj_710), .Z(n15_adj_564)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17275_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_461_i4_4_lut (.A(n2_adj_991), .B(C), .C(n7939), .D(n7943), 
         .Z(n4_adj_992)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_461_i4_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_293_i14_3_lut_4_lut (.A(n22234), .B(n7762), .C(Z_N_387[6]), 
         .D(n13_adj_940), .Z(n14_adj_877)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_293_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17269_3_lut_4_lut (.A(n22177), .B(n22091), .C(n14_adj_993), 
         .D(n10_adj_701), .Z(n15_adj_570)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17269_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_269_i14_3_lut_4_lut (.A(n22234), .B(n7762), .C(Z_N_387[0]), 
         .D(n10_adj_937), .Z(n14_adj_968)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_269_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i16467_3_lut (.A(s_2_5), .B(s_3_5), .C(instruction[4]), .Z(n19637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16467_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_361_i9_3_lut_4_lut (.A(n22101), .B(n16312), .C(n14_adj_501), 
         .D(C), .Z(n9_adj_994)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_361_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_297_i14_3_lut_4_lut (.A(n22234), .B(n7762), .C(Z_N_387[7]), 
         .D(n10_adj_926), .Z(n14_adj_597)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_297_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_108 (.A(n22304), .B(n22284), .C(n22282), 
         .D(n22307), .Z(n1[11])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_108.init = 16'h0080;
    LUT4 i16466_3_lut (.A(s_0_5), .B(s_1_5), .C(instruction[4]), .Z(n19636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16466_3_lut.init = 16'hcaca;
    LUT4 i17559_2_lut_3_lut_4_lut (.A(n22264), .B(n7876), .C(n20160), 
         .D(n7908), .Z(n19570)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17559_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 PrioSelect_489_i8_4_lut (.A(n6_adj_995), .B(n14_adj_711), .C(n7926), 
         .D(n7922), .Z(n8_adj_996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_489_i8_4_lut.init = 16'hcfca;
    LUT4 i17284_3_lut_4_lut (.A(n22183), .B(n22092), .C(n14_adj_997), 
         .D(n10_adj_998), .Z(n15_adj_552)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17284_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17528_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n7876), .C(n11714), 
         .D(n22263), .Z(n17339)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17528_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h040c;
    LUT4 i17476_2_lut_3_lut_4_lut (.A(n22264), .B(n7876), .C(n20077), 
         .D(n11714), .Z(n17362)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17476_2_lut_3_lut_4_lut.init = 16'hf0f4;
    LUT4 i17574_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n7876), .C(n7762), 
         .D(n22263), .Z(n18075)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17574_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i17563_2_lut_3_lut_4_lut (.A(n22264), .B(n7876), .C(n20164), 
         .D(n11714), .Z(n17213)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17563_2_lut_3_lut_4_lut.init = 16'hf0f4;
    LUT4 PrioSelect_309_i11_3_lut_4_lut (.A(n22235), .B(n7762), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_999)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_309_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i17566_2_lut_3_lut_4_lut (.A(n22264), .B(n7876), .C(n20167), 
         .D(n7762), .Z(n18098)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17566_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i6037_2_lut (.A(instruction[9]), .B(n8773), .Z(n8627)) /* synthesis lut_function=(!(A+!(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i6037_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_109 (.A(st_zc[1]), .B(n22283), .C(n7746), 
         .D(n22307), .Z(n1[18])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_109.init = 16'h0040;
    LUT4 i17286_3_lut_4_lut (.A(n22183), .B(n22092), .C(n14_adj_1000), 
         .D(n10_adj_1001), .Z(n15_adj_550)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17286_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n2083_bdd_4_lut_17863 (.A(n22109), .B(n2085), .C(n16312), .D(n7876), 
         .Z(n21132)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam n2083_bdd_4_lut_17863.init = 16'h1fff;
    LUT4 i17280_3_lut_4_lut (.A(n22183), .B(n22092), .C(n14_adj_1002), 
         .D(n10_adj_1003), .Z(n15_adj_556)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17280_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17290_3_lut_4_lut (.A(n22183), .B(n22092), .C(n14_adj_1004), 
         .D(n10_adj_1005), .Z(n15_adj_546)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17290_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16458_3_lut (.A(s_14_7), .B(s_15_7), .C(instruction[4]), .Z(n19628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16458_3_lut.init = 16'hcaca;
    LUT4 i16457_3_lut (.A(s_12_7), .B(s_13_7), .C(instruction[4]), .Z(n19627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16457_3_lut.init = 16'hcaca;
    LUT4 i17282_3_lut_4_lut (.A(n22183), .B(n22092), .C(n14_adj_1006), 
         .D(n10_adj_1007), .Z(n15_adj_554)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17282_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17288_3_lut_4_lut (.A(n22183), .B(n22092), .C(n14_adj_1008), 
         .D(n10_adj_1009), .Z(n15_adj_548)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17288_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_393_i9_3_lut_4_lut (.A(n22093), .B(n16312), .C(n14_adj_501), 
         .D(C), .Z(n9_adj_1010)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_393_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_493_i4_4_lut (.A(n2_adj_1011), .B(C), .C(n7940), .D(n7944), 
         .Z(n4_adj_1012)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_493_i4_4_lut.init = 16'hc0ca;
    LUT4 i17746_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n7876), .C(n16312), 
         .D(n22263), .Z(n18811)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17746_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i17304_3_lut_4_lut (.A(n22189), .B(n22094), .C(n14_adj_1013), 
         .D(n10_adj_730), .Z(n15_adj_521)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17304_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_305_i11_3_lut_4_lut (.A(n22235), .B(n7762), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1014)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_305_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i16456_3_lut (.A(s_10_7), .B(s_11_7), .C(instruction[4]), .Z(n19626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16456_3_lut.init = 16'hcaca;
    LUT4 i16455_3_lut (.A(s_8_7), .B(s_9_7), .C(instruction[4]), .Z(n19625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16455_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_525_i4_4_lut (.A(n2_adj_1015), .B(C), .C(n7941), .D(n7945), 
         .Z(n4_adj_1016)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_525_i4_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_313_i11_3_lut_4_lut (.A(n22235), .B(n7762), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1017)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_313_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i16454_3_lut (.A(s_6_7), .B(s_7_7), .C(instruction[4]), .Z(n19624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16454_3_lut.init = 16'hcaca;
    LUT4 i16453_3_lut (.A(s_4_7), .B(s_5_7), .C(instruction[4]), .Z(n19623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16453_3_lut.init = 16'hcaca;
    LUT4 i17294_3_lut_4_lut (.A(n22189), .B(n22094), .C(n14_adj_1018), 
         .D(n10_adj_719), .Z(n15_adj_537)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17294_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16452_3_lut (.A(s_2_7), .B(s_3_7), .C(instruction[4]), .Z(n19622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16452_3_lut.init = 16'hcaca;
    LUT4 i16451_3_lut (.A(s_0_7), .B(s_1_7), .C(instruction[4]), .Z(n19621)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16451_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_557_i4_4_lut (.A(n2_adj_1019), .B(C), .C(n7942), .D(n7946), 
         .Z(n4_adj_1020)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_557_i4_4_lut.init = 16'hc0ca;
    LUT4 i16443_3_lut (.A(s_14_2), .B(s_15_2), .C(instruction[4]), .Z(n19613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16443_3_lut.init = 16'hcaca;
    LUT4 i17300_3_lut_4_lut (.A(n22189), .B(n22094), .C(n14_adj_1021), 
         .D(n10_adj_728), .Z(n15_adj_525)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17300_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16442_3_lut (.A(s_12_2), .B(s_13_2), .C(instruction[4]), .Z(n19612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16442_3_lut.init = 16'hcaca;
    LUT4 i16441_3_lut (.A(s_10_2), .B(s_11_2), .C(instruction[4]), .Z(n19611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16441_3_lut.init = 16'hcaca;
    LUT4 i16440_3_lut (.A(s_8_2), .B(s_9_2), .C(instruction[4]), .Z(n19610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16440_3_lut.init = 16'hcaca;
    LUT4 i37_then_4_lut (.A(n8_adj_695), .B(instruction[16]), .C(instruction[17]), 
         .D(n8_adj_849), .Z(n22324)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C)) */ ;
    defparam i37_then_4_lut.init = 16'hfaf8;
    LUT4 i17298_3_lut_4_lut (.A(n22189), .B(n22094), .C(n14_adj_1022), 
         .D(n10_adj_727), .Z(n15_adj_533)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17298_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16439_3_lut (.A(s_6_2), .B(s_7_2), .C(instruction[4]), .Z(n19609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16439_3_lut.init = 16'hcaca;
    LUT4 i16438_3_lut (.A(s_4_2), .B(s_5_2), .C(instruction[4]), .Z(n19608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16438_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_317_i11_3_lut_4_lut (.A(n22235), .B(n7762), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1023)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_317_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_429_i16 (.BLUT(n14_adj_1024), .ALUT(n15_adj_1025), 
          .C0(n18838), .Z(n16_adj_1026)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i16437_3_lut (.A(s_2_2), .B(s_3_2), .C(instruction[4]), .Z(n19607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16437_3_lut.init = 16'hcaca;
    LUT4 i16436_3_lut (.A(s_0_2), .B(s_1_2), .C(instruction[4]), .Z(n19606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16436_3_lut.init = 16'hcaca;
    LUT4 i17302_3_lut_4_lut (.A(n22189), .B(n22094), .C(n14_adj_1027), 
         .D(n10_adj_729), .Z(n15_adj_523)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17302_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16428_3_lut (.A(s_14_4), .B(s_15_4), .C(instruction[4]), .Z(n19598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16428_3_lut.init = 16'hcaca;
    LUT4 i16427_3_lut (.A(s_12_4), .B(s_13_4), .C(instruction[4]), .Z(n19597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16427_3_lut.init = 16'hcaca;
    LUT4 i16426_3_lut (.A(s_10_4), .B(s_11_4), .C(instruction[4]), .Z(n19596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16426_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_321_i11_3_lut_4_lut (.A(n22235), .B(n7762), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1028)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_321_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i16425_3_lut (.A(s_8_4), .B(s_9_4), .C(instruction[4]), .Z(n19595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16425_3_lut.init = 16'hcaca;
    LUT4 i16424_3_lut (.A(s_6_4), .B(s_7_4), .C(instruction[4]), .Z(n19594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16424_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_325_i11_3_lut_4_lut (.A(n22235), .B(n7762), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1029)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_325_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_110 (.A(instruction[16]), .B(instruction[17]), .Z(n8070)) /* synthesis lut_function=(A+(B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[16:28])
    defparam i1_2_lut_adj_110.init = 16'heeee;
    LUT4 i16423_3_lut (.A(s_4_4), .B(s_5_4), .C(instruction[4]), .Z(n19593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16423_3_lut.init = 16'hcaca;
    LUT4 i16422_3_lut (.A(s_2_4), .B(s_3_4), .C(instruction[4]), .Z(n19592)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16422_3_lut.init = 16'hcaca;
    LUT4 i16421_3_lut (.A(s_0_4), .B(s_1_4), .C(instruction[4]), .Z(n19591)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16421_3_lut.init = 16'hcaca;
    LUT4 i16413_3_lut (.A(s_14_3), .B(s_15_3), .C(instruction[4]), .Z(n19583)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16413_3_lut.init = 16'hcaca;
    LUT4 i17602_2_lut_3_lut_4_lut (.A(n22264), .B(n7876), .C(n20203), 
         .D(n7762), .Z(n17949)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17602_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i16412_3_lut (.A(s_12_3), .B(s_13_3), .C(instruction[4]), .Z(n19582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16412_3_lut.init = 16'hcaca;
    LUT4 i16411_3_lut (.A(s_10_3), .B(s_11_3), .C(instruction[4]), .Z(n19581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16411_3_lut.init = 16'hcaca;
    LUT4 i16410_3_lut (.A(s_8_3), .B(s_9_3), .C(instruction[4]), .Z(n19580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16410_3_lut.init = 16'hcaca;
    LUT4 i17296_3_lut_4_lut (.A(n22189), .B(n22094), .C(n14_adj_1030), 
         .D(n10_adj_720), .Z(n15_adj_535)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17296_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16409_3_lut (.A(s_6_3), .B(s_7_3), .C(instruction[4]), .Z(n19579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16409_3_lut.init = 16'hcaca;
    LUT4 i16408_3_lut (.A(s_4_3), .B(s_5_3), .C(instruction[4]), .Z(n19578)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16408_3_lut.init = 16'hcaca;
    LUT4 i16407_3_lut (.A(s_2_3), .B(s_3_3), .C(instruction[4]), .Z(n19577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16407_3_lut.init = 16'hcaca;
    LUT4 i16406_3_lut (.A(s_0_3), .B(s_1_3), .C(instruction[4]), .Z(n19576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16406_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_425_i9_3_lut_4_lut (.A(n22095), .B(n16312), .C(n14_adj_501), 
         .D(C), .Z(n9_adj_1031)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_425_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i17317_3_lut_4_lut (.A(n22195), .B(n22096), .C(n14_adj_1032), 
         .D(n10_adj_1033), .Z(n15_adj_498)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17317_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17307_3_lut_4_lut (.A(n22195), .B(n22096), .C(n14_adj_1034), 
         .D(n10_adj_1035), .Z(n15_adj_510)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17307_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_329_i11_3_lut_4_lut (.A(n22236), .B(n7762), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1036)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_329_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 n2083_bdd_4_lut_17800 (.A(n22109), .B(n2085), .C(n11714), .D(n7726), 
         .Z(n20914)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam n2083_bdd_4_lut_17800.init = 16'hf1ff;
    LUT4 i17313_3_lut_4_lut (.A(n22195), .B(n22096), .C(n14_adj_1037), 
         .D(n10_adj_1038), .Z(n15_adj_504)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17313_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n10_bdd_4_lut (.A(n10_adj_812), .B(instruction[15]), .C(instruction[16]), 
         .D(instruction[17]), .Z(n21529)) /* synthesis lut_function=(A (B (D)+!B (C+!(D)))) */ ;
    defparam n10_bdd_4_lut.init = 16'ha822;
    LUT4 i37_else_4_lut (.A(n8050), .B(n8_adj_695), .C(instruction[16]), 
         .D(instruction[17]), .Z(n22323)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i37_else_4_lut.init = 16'hfff8;
    LUT4 i1_4_lut (.A(n24), .B(n21187), .C(n4_adj_1039), .D(n4_adj_1040), 
         .Z(n63_adj_1041)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfcec;
    LUT4 i1562_3_lut_4_lut (.A(n8627), .B(n11714), .C(n7_adj_473), .D(n7_adj_609), 
         .Z(n10_adj_1042)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1562_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_827_8 (.A0(instruction[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(instruction[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14285), .COUT(n14286), .S0(C_N_342[6]), 
          .S1(C_N_342[7]));   // f:/home/mini-mcu/step_fpga/mcu.v(281[97:106])
    defparam add_827_8.INIT0 = 16'hfaaa;
    defparam add_827_8.INIT1 = 16'hfaaa;
    defparam add_827_8.INJECT1_0 = "NO";
    defparam add_827_8.INJECT1_1 = "NO";
    LUT4 i17311_3_lut_4_lut (.A(n22195), .B(n22096), .C(n14_adj_1043), 
         .D(n10_adj_1044), .Z(n15_adj_506)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17311_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17315_3_lut_4_lut (.A(n22195), .B(n22096), .C(n14_adj_1045), 
         .D(n10_adj_1046), .Z(n15_adj_502)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17315_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17309_3_lut_4_lut (.A(n22195), .B(n22096), .C(n14_adj_1047), 
         .D(n10_adj_1048), .Z(n15_adj_508)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17309_3_lut_4_lut.init = 16'hf1e0;
    CCU2D add_827_6 (.A0(instruction[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(instruction[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14284), .COUT(n14285), .S0(C_N_342[4]), 
          .S1(C_N_342[5]));   // f:/home/mini-mcu/step_fpga/mcu.v(281[97:106])
    defparam add_827_6.INIT0 = 16'hfaaa;
    defparam add_827_6.INIT1 = 16'hfaaa;
    defparam add_827_6.INJECT1_0 = "NO";
    defparam add_827_6.INJECT1_1 = "NO";
    LUT4 PrioSelect_301_i11_3_lut_4_lut (.A(n22236), .B(n7762), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1049)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_301_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_457_i9_3_lut_4_lut (.A(n22097), .B(n16312), .C(n14_adj_501), 
         .D(C), .Z(n9_adj_1050)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_457_i9_3_lut_4_lut.init = 16'hf780;
    CCU2D add_827_4 (.A0(instruction[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(instruction[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14283), .COUT(n14284), .S0(C_N_342[2]), 
          .S1(C_N_342[3]));   // f:/home/mini-mcu/step_fpga/mcu.v(281[97:106])
    defparam add_827_4.INIT0 = 16'hfaaa;
    defparam add_827_4.INIT1 = 16'hfaaa;
    defparam add_827_4.INJECT1_0 = "NO";
    defparam add_827_4.INJECT1_1 = "NO";
    LUT4 i17723_2_lut_3_lut_4_lut (.A(n22264), .B(n7876), .C(n20324), 
         .D(n16312), .Z(n18834)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17723_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i17331_3_lut_4_lut (.A(n22213), .B(n22098), .C(n14_adj_1051), 
         .D(n10_adj_749), .Z(n15_adj_466)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17331_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6096_2_lut_3_lut_4_lut (.A(n160), .B(instruction[3]), .C(n7646), 
         .D(instruction[8]), .Z(n8773)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i6096_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i17573_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22237), .B(n7762), .C(n22235), 
         .D(n22236), .Z(n18090)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17573_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hccc8;
    LUT4 PrioSelect_301_i12_3_lut_4_lut (.A(n22237), .B(n7762), .C(Z_N_378[0]), 
         .D(n11_adj_1049), .Z(n12_adj_1052)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_301_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17321_3_lut_4_lut (.A(n22213), .B(n22098), .C(n14_adj_1053), 
         .D(n10_adj_738), .Z(n15_adj_483)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17321_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_329_i12_3_lut_4_lut (.A(n22237), .B(n7762), .C(Z_N_378[7]), 
         .D(n11_adj_1036), .Z(n12_adj_578)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_329_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17757_2_lut_3_lut_4_lut (.A(n22264), .B(n7876), .C(n20358), 
         .D(n16312), .Z(n18685)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17757_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i17567_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n7876), .C(n7908), 
         .D(n22263), .Z(n19547)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17567_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i17327_3_lut_4_lut (.A(n22213), .B(n22098), .C(n14_adj_1054), 
         .D(n10_adj_745), .Z(n15_adj_471)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17327_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6013_2_lut_rep_552_3_lut_4_lut (.A(n160), .B(instruction[3]), 
         .C(n7646), .D(n7726), .Z(n22119)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i6013_2_lut_rep_552_3_lut_4_lut.init = 16'h8000;
    LUT4 i17531_2_lut_rep_519_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n7876), 
         .C(n11714), .D(n22268), .Z(n22086)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17531_2_lut_rep_519_3_lut_3_lut_4_lut_4_lut.init = 16'h040c;
    LUT4 i17325_3_lut_4_lut (.A(n22213), .B(n22098), .C(n14_adj_1055), 
         .D(n10_adj_741), .Z(n15_adj_474)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17325_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17577_2_lut_rep_523_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n7876), 
         .C(n7762), .D(n22268), .Z(n22090)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17577_2_lut_rep_523_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i17329_3_lut_4_lut (.A(n22213), .B(n22098), .C(n14_adj_1056), 
         .D(n10_adj_747), .Z(n15_adj_469)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17329_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_then_3_lut (.A(instruction[17]), .B(instruction[14]), 
         .C(instruction[15]), .Z(n22327)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_4_lut_then_3_lut.init = 16'h8080;
    LUT4 i17323_3_lut_4_lut (.A(n22213), .B(n22098), .C(n14_adj_1057), 
         .D(n10_adj_740), .Z(n15_adj_477)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17323_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17358_3_lut_4_lut (.A(n22122), .B(n22099), .C(n14_adj_1058), 
         .D(n10_adj_1059), .Z(n15_adj_1060)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17358_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17348_3_lut_4_lut (.A(n22122), .B(n22099), .C(n14_adj_1061), 
         .D(n10_adj_1062), .Z(n15_adj_1063)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17348_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_305_i12_3_lut_4_lut (.A(n22238), .B(n7762), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1064)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_305_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_309_i12_3_lut_4_lut (.A(n22238), .B(n7762), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1065)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_309_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17749_2_lut_rep_529_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n7876), 
         .C(n16312), .D(n22268), .Z(n22096)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17749_2_lut_rep_529_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 PrioSelect_313_i12_3_lut_4_lut (.A(n22238), .B(n7762), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1066)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_313_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17570_2_lut_rep_533_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n7876), 
         .C(n7908), .D(n22268), .Z(n22100)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17570_2_lut_rep_533_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i17354_3_lut_4_lut (.A(n22122), .B(n22099), .C(n14_adj_1067), 
         .D(n10_adj_1068), .Z(n15_adj_1069)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17354_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i8805_4_lut_then_3_lut (.A(n8_adj_695), .B(instruction[17]), .C(instruction[15]), 
         .Z(n22309)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i8805_4_lut_then_3_lut.init = 16'hefef;
    LUT4 PrioSelect_317_i12_3_lut_4_lut (.A(n22238), .B(n7762), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1070)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_317_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i8544_4_lut (.A(s_15_0), .B(n9), .C(n9_adj_1), .D(n7908), .Z(n2_adj_1019)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8544_4_lut.init = 16'hceaa;
    LUT4 i1_3_lut_4_lut_else_3_lut (.A(instruction[17]), .B(instruction[14]), 
         .C(instruction[15]), .D(instruction[13]), .Z(n22326)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)))+!A (B+(D)))) */ ;
    defparam i1_3_lut_4_lut_else_3_lut.init = 16'h02b3;
    LUT4 i3178_3_lut_4_lut (.A(n22227), .B(n22281), .C(n13_adj_739), .D(n13_adj_731), 
         .Z(n10_adj_1073)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i3178_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_321_i12_3_lut_4_lut (.A(n22238), .B(n7762), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1074)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_321_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_325_i12_3_lut_4_lut (.A(n22238), .B(n7762), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1075)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_325_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17352_3_lut_4_lut (.A(n22122), .B(n22099), .C(n14_adj_1076), 
         .D(n10_adj_1077), .Z(n15_adj_1078)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17352_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17356_3_lut_4_lut (.A(n22122), .B(n22099), .C(n14_adj_1079), 
         .D(n10_adj_1080), .Z(n15_adj_1081)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17356_3_lut_4_lut.init = 16'hf1e0;
    PFUMX PrioSelect_365_i16 (.BLUT(n14_adj_1082), .ALUT(n15_adj_1083), 
          .C0(n18321), .Z(n16_adj_1084)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17350_3_lut_4_lut (.A(n22122), .B(n22099), .C(n14_adj_1085), 
         .D(n10_adj_1086), .Z(n15_adj_1087)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17350_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17372_3_lut_4_lut (.A(n22116), .B(n22100), .C(n14_adj_1088), 
         .D(n10_adj_1089), .Z(n15_adj_1090)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17372_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_301_i15_3_lut_4_lut (.A(n22238), .B(n7762), .C(n1108[0]), 
         .D(n5_adj_1091), .Z(n15_adj_1092)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_301_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i17362_3_lut_4_lut (.A(n22116), .B(n22100), .C(n14_adj_1093), 
         .D(n10_adj_1094), .Z(n15_adj_1095)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17362_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_329_i15_3_lut_4_lut (.A(n22238), .B(n7762), .C(n1108[7]), 
         .D(n9_adj_956), .Z(n15_adj_575)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_329_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i3194_3_lut_4_lut (.A(n22227), .B(n22281), .C(n13_adj_516), .D(n13_adj_736), 
         .Z(n10_adj_1096)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i3194_3_lut_4_lut.init = 16'hf780;
    LUT4 i3210_3_lut_4_lut (.A(n22227), .B(n22281), .C(n13_adj_744), .D(n13_adj_739), 
         .Z(n10_adj_1097)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i3210_3_lut_4_lut.init = 16'hf780;
    LUT4 i17368_3_lut_4_lut (.A(n22116), .B(n22100), .C(n14_adj_1098), 
         .D(n10_adj_1097), .Z(n15_adj_1099)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17368_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_329_i10_3_lut_4_lut (.A(n22239), .B(n7762), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1100)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_329_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i17366_3_lut_4_lut (.A(n22116), .B(n22100), .C(n14_adj_1101), 
         .D(n10_adj_1096), .Z(n15_adj_1102)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17366_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_561_i17_3_lut_4_lut (.A(n22266), .B(n22281), .C(in_port[1]), 
         .D(n16_adj_1103), .Z(n17_adj_1104)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_561_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17370_3_lut_4_lut (.A(n22116), .B(n22100), .C(n14_adj_1105), 
         .D(n10_adj_517), .Z(n15_adj_1106)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17370_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n2083_bdd_4_lut_17816 (.A(n22109), .B(n2085), .C(n11714), .D(n16392), 
         .Z(n20955)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam n2083_bdd_4_lut_17816.init = 16'hf1ff;
    LUT4 i2250_3_lut_4_lut (.A(n22239), .B(n7762), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1107)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i2250_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_565_i17_3_lut_4_lut (.A(n22266), .B(n22281), .C(in_port[2]), 
         .D(n16_adj_1108), .Z(n17_adj_1109)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_565_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17364_3_lut_4_lut (.A(n22116), .B(n22100), .C(n14_adj_1110), 
         .D(n10_adj_1073), .Z(n15_adj_1111)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17364_3_lut_4_lut.init = 16'hf1e0;
    LUT4 PrioSelect_569_i17_3_lut_4_lut (.A(n22266), .B(n22281), .C(in_port[3]), 
         .D(n16_adj_1112), .Z(n17_adj_1113)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_569_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_573_i17_3_lut_4_lut (.A(n22266), .B(n22281), .C(in_port[4]), 
         .D(n16_adj_1114), .Z(n17_adj_1115)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_573_i17_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_827_2 (.A0(C), .B0(instruction[0]), .C0(GND_net), .D0(GND_net), 
          .A1(instruction[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n14283), .S1(C_N_342[1]));   // f:/home/mini-mcu/step_fpga/mcu.v(281[97:106])
    defparam add_827_2.INIT0 = 16'h7000;
    defparam add_827_2.INIT1 = 16'hfaaa;
    defparam add_827_2.INJECT1_0 = "NO";
    defparam add_827_2.INJECT1_1 = "NO";
    LUT4 PrioSelect_489_i9_3_lut_4_lut (.A(n22101), .B(n7908), .C(n14_adj_501), 
         .D(C), .Z(n9_adj_1116)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_489_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_577_i17_3_lut_4_lut (.A(n22266), .B(n22281), .C(in_port[5]), 
         .D(n16_adj_1117), .Z(n17_adj_1118)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_577_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 n2083_bdd_4_lut_17883 (.A(n22109), .B(n2085), .C(n7908), .D(n11778), 
         .Z(n21170)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;
    defparam n2083_bdd_4_lut_17883.init = 16'hff1f;
    CCU2D add_632_5 (.A0(instruction[3]), .B0(n7_c), .C0(instruction[11]), 
          .D0(n14), .A1(instruction[4]), .B1(n7_adj_462), .C1(instruction[11]), 
          .D1(n14_adj_463), .CIN(n14262), .COUT(n14263), .S0(Z_N_367[3]), 
          .S1(Z_N_367[4]));   // f:/home/mini-mcu/step_fpga/mcu.v(263[59:70])
    defparam add_632_5.INIT0 = 16'h56a6;
    defparam add_632_5.INIT1 = 16'h56a6;
    defparam add_632_5.INJECT1_0 = "NO";
    defparam add_632_5.INJECT1_1 = "NO";
    LUT4 PrioSelect_581_i17_3_lut_4_lut (.A(n22266), .B(n22281), .C(in_port[6]), 
         .D(n16_adj_1119), .Z(n17_adj_1120)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_581_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i14200_3_lut_3_lut_4_lut (.A(n2075), .B(n11778), .C(n8627), .D(n7762), 
         .Z(n17370)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(223[39:43])
    defparam i14200_3_lut_3_lut_4_lut.init = 16'h0dff;
    LUT4 i14936_3_lut_3_lut_4_lut (.A(n2075), .B(n11778), .C(n16312), 
         .D(n8627), .Z(n18106)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(223[39:43])
    defparam i14936_3_lut_3_lut_4_lut.init = 16'h0fdf;
    LUT4 PrioSelect_325_i13_3_lut_4_lut (.A(n22239), .B(n7762), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1121)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_325_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i8535_4_lut (.A(s_14_0), .B(n7), .C(n7_adj_2), .D(n7908), .Z(n2_adj_1015)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8535_4_lut.init = 16'hceaa;
    LUT4 i15672_3_lut_3_lut_4_lut (.A(n2075), .B(n11778), .C(n7908), .D(n8627), 
         .Z(n18842)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(223[39:43])
    defparam i15672_3_lut_3_lut_4_lut.init = 16'h0fdf;
    LUT4 instruction_13__bdd_4_lut (.A(instruction[14]), .B(instruction[12]), 
         .C(instruction[15]), .D(instruction[16]), .Z(n21186)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam instruction_13__bdd_4_lut.init = 16'hc2c0;
    LUT4 PrioSelect_321_i13_3_lut_4_lut (.A(n22239), .B(n7762), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1124)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_321_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_317_i13_3_lut_4_lut (.A(n22239), .B(n7762), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1125)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_317_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i17666_4_lut (.A(n22214), .B(n22219), .C(n22218), .D(n19164), 
         .Z(n20268)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17666_4_lut.init = 16'habaa;
    LUT4 i8524_4_lut (.A(s_13_0), .B(n10), .C(n10_adj_3), .D(n7908), 
         .Z(n2_adj_1011)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8524_4_lut.init = 16'hceaa;
    LUT4 PrioSelect_313_i13_3_lut_4_lut (.A(n22239), .B(n7762), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1128)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_313_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i17748_2_lut_3_lut_4_lut (.A(n16312), .B(n22266), .C(n20349), 
         .D(n7876), .Z(n18809)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;
    defparam i17748_2_lut_3_lut_4_lut.init = 16'hf2f0;
    LUT4 PrioSelect_309_i13_3_lut_4_lut (.A(n22239), .B(n7762), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1129)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_309_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i15974_4_lut (.A(n22217), .B(n22216), .C(n22215), .D(n213[13]), 
         .Z(n19164)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15974_4_lut.init = 16'h5554;
    LUT4 PrioSelect_305_i13_3_lut_4_lut (.A(n22239), .B(n7762), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1130)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_305_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i17765_2_lut_3_lut_4_lut (.A(n16312), .B(n22266), .C(n20366), 
         .D(n16392), .Z(n18625)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;
    defparam i17765_2_lut_3_lut_4_lut.init = 16'hf2f0;
    PFUMX PrioSelect_301_i16 (.BLUT(n14_adj_1131), .ALUT(n15_adj_1092), 
          .C0(n18102), .Z(n16_adj_1132)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i13832_3_lut_3_lut_4_lut (.A(n2075), .B(n16392), .C(n11714), 
         .D(n8647), .Z(n17002)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C+!(D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(223[39:43])
    defparam i13832_3_lut_3_lut_4_lut.init = 16'hf0f7;
    LUT4 i14568_3_lut_3_lut_4_lut (.A(n2075), .B(n16392), .C(n8647), .D(n7762), 
         .Z(n17738)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(223[39:43])
    defparam i14568_3_lut_3_lut_4_lut.init = 16'h07ff;
    LUT4 i15304_3_lut_3_lut_4_lut (.A(n2075), .B(n16392), .C(n16312), 
         .D(n8647), .Z(n18474)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(223[39:43])
    defparam i15304_3_lut_3_lut_4_lut.init = 16'h0f7f;
    LUT4 i3162_3_lut_4_lut (.A(n22227), .B(n22281), .C(n13_adj_736), .D(n5_adj_737), 
         .Z(n10_adj_1094)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i3162_3_lut_4_lut.init = 16'hf780;
    LUT4 i8521_4_lut (.A(s_12_7), .B(n7931), .C(n13_adj_515), .D(n6886), 
         .Z(n6_adj_995)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8521_4_lut.init = 16'h3022;
    LUT4 PrioSelect_305_i14_3_lut_4_lut (.A(n22240), .B(n7762), .C(Z_N_387[1]), 
         .D(n13_adj_1130), .Z(n14_adj_910)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_305_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_309_i14_3_lut_4_lut (.A(n22240), .B(n7762), .C(Z_N_387[2]), 
         .D(n13_adj_1129), .Z(n14_adj_931)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_309_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_313_i14_3_lut_4_lut (.A(n22240), .B(n7762), .C(Z_N_387[3]), 
         .D(n13_adj_1128), .Z(n14_adj_920)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_313_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_317_i14_3_lut_4_lut (.A(n22240), .B(n7762), .C(Z_N_387[4]), 
         .D(n13_adj_1125), .Z(n14_adj_912)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_317_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_321_i14_3_lut_4_lut (.A(n22240), .B(n7762), .C(Z_N_387[5]), 
         .D(n13_adj_1124), .Z(n14_adj_929)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_321_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17488_2_lut_3_lut_4_lut (.A(n16312), .B(n22266), .C(n20089), 
         .D(n7726), .Z(n18361)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;
    defparam i17488_2_lut_3_lut_4_lut.init = 16'hf2f0;
    CCU2D add_21_3 (.A0(address[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(address[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14265), .COUT(n14266), .S0(n18[1]), .S1(n18[2]));   // f:/home/mini-mcu/step_fpga/mcu.v(217[27:35])
    defparam add_21_3.INIT0 = 16'h5aaa;
    defparam add_21_3.INIT1 = 16'h5aaa;
    defparam add_21_3.INJECT1_0 = "NO";
    defparam add_21_3.INJECT1_1 = "NO";
    LUT4 PrioSelect_325_i14_3_lut_4_lut (.A(n22240), .B(n7762), .C(Z_N_387[6]), 
         .D(n13_adj_1121), .Z(n14_adj_906)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_325_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_301_i14_3_lut_4_lut (.A(n22240), .B(n7762), .C(Z_N_387[0]), 
         .D(n10_adj_1107), .Z(n14_adj_1131)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_301_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i16040_3_lut_4_lut (.A(n2075), .B(n16392), .C(n7908), .D(n22083), 
         .Z(n19210)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(223[39:43])
    defparam i16040_3_lut_4_lut.init = 16'h007f;
    LUT4 n21795_bdd_2_lut_4_lut (.A(s_N_294[3]), .B(n10_adj_1133), .C(s_N_294[6]), 
         .D(n21795), .Z(n21796)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(227[81:100])
    defparam n21795_bdd_2_lut_4_lut.init = 16'h0100;
    LUT4 PrioSelect_329_i14_3_lut_4_lut (.A(n22240), .B(n7762), .C(Z_N_387[7]), 
         .D(n10_adj_1100), .Z(n14_adj_574)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_329_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i8805_4_lut_else_3_lut (.A(n8_adj_849), .B(n8_adj_695), .C(instruction[17]), 
         .D(instruction[15]), .Z(n22308)) /* synthesis lut_function=(A (B+(C))+!A (B (C+!(D))+!B (C))) */ ;
    defparam i8805_4_lut_else_3_lut.init = 16'hf8fc;
    LUT4 n21186_bdd_2_lut (.A(n21186), .B(instruction[13]), .Z(n21187)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n21186_bdd_2_lut.init = 16'h2222;
    LUT4 i8514_4_lut (.A(s_12_0), .B(n8), .C(n8_adj_4), .D(n7908), .Z(n2_adj_991)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8514_4_lut.init = 16'hceaa;
    LUT4 PrioSelect_341_i11_3_lut_4_lut (.A(n22245), .B(n16312), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1136)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_341_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17543_2_lut_3_lut_4_lut (.A(n16312), .B(n22266), .C(n20144), 
         .D(n11778), .Z(n18257)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;
    defparam i17543_2_lut_3_lut_4_lut.init = 16'hf0f2;
    LUT4 PrioSelect_337_i11_3_lut_4_lut (.A(n22245), .B(n16312), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1137)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_337_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i6023_2_lut_rep_551_3_lut_4_lut (.A(n160), .B(instruction[3]), 
         .C(n7646), .D(n7876), .Z(n22118)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i6023_2_lut_rep_551_3_lut_4_lut.init = 16'h8000;
    LUT4 PrioSelect_345_i11_3_lut_4_lut (.A(n22245), .B(n16312), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1138)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_345_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_349_i11_3_lut_4_lut (.A(n22245), .B(n16312), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1139)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_349_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8505_4_lut (.A(s_11_0), .B(n9), .C(n9_adj_1), .D(n16312), 
         .Z(n2_adj_971)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8505_4_lut.init = 16'hceaa;
    LUT4 PrioSelect_353_i11_3_lut_4_lut (.A(n22245), .B(n16312), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1140)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_353_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_4_lut_4_lut (.A(n22261), .B(n11778), .C(n7908), .D(n22205), 
         .Z(clk_in_c_enable_88)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+((D)+!C)))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h2030;
    LUT4 i14016_3_lut_4_lut_4_lut_4_lut (.A(n7876), .B(n22227), .C(n2075), 
         .D(n11714), .Z(n17186)) /* synthesis lut_function=((B (D)+!B ((D)+!C))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14016_3_lut_4_lut_4_lut_4_lut.init = 16'hff57;
    LUT4 PrioSelect_357_i11_3_lut_4_lut (.A(n22245), .B(n16312), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1141)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_357_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8502_4_lut (.A(s_10_7), .B(n16330), .C(n14_adj_709), .D(n16356), 
         .Z(n6_adj_958)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8502_4_lut.init = 16'h3022;
    LUT4 i1_2_lut_4_lut_4_lut_adj_111 (.A(n22261), .B(n11778), .C(n7762), 
         .D(n22205), .Z(clk_in_c_enable_40)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+((D)+!C)))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_111.init = 16'h2030;
    LUT4 i1_4_lut_4_lut_adj_112 (.A(n22261), .B(n11778), .C(n22205), .D(n16312), 
         .Z(clk_in_c_enable_64)) /* synthesis lut_function=(!(A (B+!(D))+!A (B+(C+!(D))))) */ ;
    defparam i1_4_lut_4_lut_adj_112.init = 16'h2300;
    LUT4 i16224_3_lut_4_lut (.A(n2075), .B(n7876), .C(n7908), .D(n22117), 
         .Z(n19394)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(223[39:43])
    defparam i16224_3_lut_4_lut.init = 16'h007f;
    PFUMX PrioSelect_237_i16 (.BLUT(n14_adj_734), .ALUT(n15_adj_1142), .C0(n17734), 
          .Z(n16_adj_1143)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_361_i11_3_lut_4_lut (.A(n22246), .B(n16312), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1144)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_361_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_333_i11_3_lut_4_lut (.A(n22246), .B(n16312), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1145)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_333_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17576_2_lut_3_lut_4_lut (.A(n7762), .B(n22266), .C(n20177), 
         .D(n7876), .Z(n18073)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;
    defparam i17576_2_lut_3_lut_4_lut.init = 16'hf2f0;
    LUT4 i14752_3_lut_4_lut_4_lut_4_lut (.A(n7876), .B(n22227), .C(n2075), 
         .D(n7762), .Z(n17922)) /* synthesis lut_function=(!(A (B (D)+!B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14752_3_lut_4_lut_4_lut_4_lut.init = 16'h57ff;
    LUT4 i15488_3_lut_4_lut_4_lut_4_lut (.A(n7876), .B(n22227), .C(n2075), 
         .D(n16312), .Z(n18658)) /* synthesis lut_function=(!(A (B (D)+!B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15488_3_lut_4_lut_4_lut_4_lut.init = 16'h57ff;
    LUT4 i17534_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22248), .B(n16312), .C(n22245), 
         .D(n22246), .Z(n18274)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17534_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h4ccc;
    LUT4 i8496_4_lut (.A(s_10_0), .B(n7), .C(n7_adj_2), .D(n16312), 
         .Z(n2_adj_949)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8496_4_lut.init = 16'hceaa;
    LUT4 PrioSelect_361_i12_3_lut_4_lut (.A(n22248), .B(n16312), .C(Z_N_378[7]), 
         .D(n11_adj_1144), .Z(n12_adj_1146)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_361_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_333_i12_3_lut_4_lut (.A(n22248), .B(n16312), .C(Z_N_378[0]), 
         .D(n11_adj_1145), .Z(n12_adj_1147)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_333_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8487_4_lut (.A(s_9_0), .B(n10), .C(n10_adj_3), .D(n16312), 
         .Z(n2_adj_947)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8487_4_lut.init = 16'hceaa;
    LUT4 PrioSelect_109_i5_3_lut_4_lut (.A(n22119), .B(n11714), .C(n7_adj_479), 
         .D(n7_adj_473), .Z(n5_adj_1148)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_109_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut_4_lut_adj_113 (.A(st_zc[1]), .B(n22283), .C(n22282), 
         .D(n22307), .Z(n1[14])) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_113.init = 16'h4000;
    CCU2D add_21_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(address[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n14265), .S1(n18[0]));   // f:/home/mini-mcu/step_fpga/mcu.v(217[27:35])
    defparam add_21_1.INIT0 = 16'hF000;
    defparam add_21_1.INIT1 = 16'h5555;
    defparam add_21_1.INJECT1_0 = "NO";
    defparam add_21_1.INJECT1_1 = "NO";
    LUT4 PrioSelect_337_i12_3_lut_4_lut (.A(n22250), .B(n16312), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1149)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_337_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13648_3_lut_4_lut_4_lut_4_lut (.A(n7726), .B(n22227), .C(n2075), 
         .D(n11714), .Z(n16818)) /* synthesis lut_function=((B (D)+!B ((D)+!C))+!A) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i13648_3_lut_4_lut_4_lut_4_lut.init = 16'hff57;
    LUT4 i8567_4_lut (.A(n22313), .B(rst_n_in), .C(st[3]), .D(n1124), 
         .Z(n3[3])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam i8567_4_lut.init = 16'hc088;
    LUT4 i17657_2_lut_3_lut_4_lut (.A(n7762), .B(n22266), .C(n20258), 
         .D(n16392), .Z(n17889)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;
    defparam i17657_2_lut_3_lut_4_lut.init = 16'hf2f0;
    LUT4 i2_4_lut_adj_114 (.A(n16122), .B(n206), .C(n103), .D(instruction[0]), 
         .Z(n16123)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[26:31])
    defparam i2_4_lut_adj_114.init = 16'hfbfa;
    LUT4 PrioSelect_341_i12_3_lut_4_lut (.A(n22250), .B(n16312), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1150)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_341_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_345_i12_3_lut_4_lut (.A(n22250), .B(n16312), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1151)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_345_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8484_4_lut (.A(s_8_7), .B(n16336), .C(n14_adj_709), .D(n16354), 
         .Z(n6_adj_945)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8484_4_lut.init = 16'h3022;
    LUT4 i17711_2_lut_3_lut_4_lut (.A(n7762), .B(n22266), .C(n20312), 
         .D(n7726), .Z(n17705)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;
    defparam i17711_2_lut_3_lut_4_lut.init = 16'hf2f0;
    LUT4 PrioSelect_349_i12_3_lut_4_lut (.A(n22250), .B(n16312), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1152)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_349_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1594_3_lut_4_lut (.A(n22119), .B(n11714), .C(n7_adj_481), .D(n7_adj_500), 
         .Z(n10_adj_758)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1594_3_lut_4_lut.init = 16'hfd20;
    LUT4 i14384_3_lut_4_lut_4_lut_4_lut (.A(n7726), .B(n22227), .C(n2075), 
         .D(n7762), .Z(n17554)) /* synthesis lut_function=(!(A (B (D)+!B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14384_3_lut_4_lut_4_lut_4_lut.init = 16'h57ff;
    LUT4 i17770_2_lut_3_lut_4_lut (.A(n7762), .B(n22266), .C(n20371), 
         .D(n11778), .Z(n17521)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;
    defparam i17770_2_lut_3_lut_4_lut.init = 16'hf0f2;
    LUT4 PrioSelect_353_i12_3_lut_4_lut (.A(n22250), .B(n16312), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1153)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_353_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_357_i12_3_lut_4_lut (.A(n22250), .B(n16312), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1154)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_357_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i15120_3_lut_4_lut_4_lut_4_lut (.A(n7726), .B(n22227), .C(n2075), 
         .D(n16312), .Z(n18290)) /* synthesis lut_function=(!(A (B (D)+!B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15120_3_lut_4_lut_4_lut_4_lut.init = 16'h57ff;
    LUT4 i15856_3_lut_4_lut_4_lut_4_lut (.A(n7726), .B(n22227), .C(n2075), 
         .D(n7908), .Z(n19026)) /* synthesis lut_function=(!(A (B (D)+!B (C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15856_3_lut_4_lut_4_lut_4_lut.init = 16'h57ff;
    LUT4 mux_308_i1_3_lut (.A(n18[0]), .B(instruction[0]), .C(n1339), 
         .Z(n1194[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i1_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_333_i15_3_lut_4_lut (.A(n22250), .B(n16312), .C(n1108[0]), 
         .D(n5_adj_1155), .Z(n15_adj_966)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_333_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8185_4_lut (.A(n2324), .B(rst_n_in), .C(n2325), .D(n2323), 
         .Z(n1742[0])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8185_4_lut.init = 16'hc088;
    LUT4 PrioSelect_361_i15_3_lut_4_lut (.A(n22250), .B(n16312), .C(n1108[7]), 
         .D(n9_adj_994), .Z(n15_adj_559)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_361_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1610_3_lut_4_lut (.A(n22119), .B(n11714), .C(n7_c), .D(n7_adj_479), 
         .Z(n10_adj_774)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1610_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_308_i12_3_lut (.A(n18[11]), .B(instruction[11]), .C(n1339), 
         .Z(n1194[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i12_3_lut.init = 16'hcaca;
    CCU2D add_632_9 (.A0(instruction[7]), .B0(n7_adj_473), .C0(instruction[11]), 
          .D0(n14_adj_711), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14264), .S0(Z_N_367[7]), .S1(C_N_338[8]));   // f:/home/mini-mcu/step_fpga/mcu.v(263[59:70])
    defparam add_632_9.INIT0 = 16'h56a6;
    defparam add_632_9.INIT1 = 16'h0000;
    defparam add_632_9.INJECT1_0 = "NO";
    defparam add_632_9.INJECT1_1 = "NO";
    LUT4 i8478_4_lut (.A(s_8_0), .B(n8), .C(n8_adj_4), .D(n16312), .Z(n2_adj_941)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8478_4_lut.init = 16'hceaa;
    LUT4 i8564_4_lut (.A(n2346), .B(rst_n_in), .C(n2347), .D(n2323), 
         .Z(n1742[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8564_4_lut.init = 16'hc088;
    LUT4 i1626_3_lut_4_lut (.A(n22119), .B(n11714), .C(n7_adj_462), .D(n7_adj_481), 
         .Z(n10_adj_768)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1626_3_lut_4_lut.init = 16'hfd20;
    LUT4 i4_4_lut (.A(n7_adj_837), .B(clk_in_c_enable_174), .C(instruction[12]), 
         .D(n20074), .Z(n14459)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i4_4_lut.init = 16'hbfff;
    LUT4 i1_2_lut_3_lut_4_lut_adj_115 (.A(st_zc[1]), .B(n22283), .C(n22285), 
         .D(n22307), .Z(n1[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_115.init = 16'h0400;
    LUT4 mux_308_i11_3_lut (.A(n18[10]), .B(instruction[10]), .C(n1339), 
         .Z(n1194[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i11_3_lut.init = 16'hcaca;
    LUT4 i1642_3_lut_4_lut (.A(n22119), .B(n11714), .C(n7_adj_609), .D(n7_c), 
         .Z(n10_adj_761)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1642_3_lut_4_lut.init = 16'hfd20;
    LUT4 i8563_4_lut (.A(n2344), .B(rst_n_in), .C(n2345), .D(n2323), 
         .Z(n1742[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8563_4_lut.init = 16'hc088;
    LUT4 mux_308_i10_3_lut (.A(n18[9]), .B(instruction[9]), .C(n1339), 
         .Z(n1194[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i10_3_lut.init = 16'hcaca;
    LUT4 i8562_4_lut (.A(n2342), .B(rst_n_in), .C(n2343), .D(n2323), 
         .Z(n1742[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8562_4_lut.init = 16'hc088;
    LUT4 PrioSelect_361_i10_3_lut_4_lut (.A(n22252), .B(n16312), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1156)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_361_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1658_3_lut_4_lut (.A(n22119), .B(n11714), .C(n7_adj_476), .D(n7_adj_462), 
         .Z(n10_adj_771)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1658_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2362_3_lut_4_lut (.A(n22252), .B(n16312), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1157)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i2362_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8469_4_lut (.A(s_7_0), .B(n9), .C(n9_adj_1), .D(n7762), .Z(n2_adj_938)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8469_4_lut.init = 16'hceaa;
    LUT4 i1674_3_lut_4_lut (.A(n22119), .B(n11714), .C(n7_adj_473), .D(n7_adj_609), 
         .Z(n10_adj_751)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1674_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_529_i12_3_lut_4_lut (.A(n22232), .B(n7908), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1158)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_529_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_173_i5_3_lut_4_lut (.A(n22118), .B(n11714), .C(n7_adj_479), 
         .D(n7_adj_473), .Z(n5_adj_1159)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_173_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_357_i13_3_lut_4_lut (.A(n22252), .B(n16312), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1160)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_357_i13_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_173_i16 (.BLUT(n14_adj_1161), .ALUT(n15_adj_1162), 
          .C0(n17366), .Z(n16_adj_1163)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_533_i12_3_lut_4_lut (.A(n22232), .B(n7908), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1164)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_533_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_537_i12_3_lut_4_lut (.A(n22232), .B(n7908), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1165)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_537_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_353_i13_3_lut_4_lut (.A(n22252), .B(n16312), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1166)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_353_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_349_i13_3_lut_4_lut (.A(n22252), .B(n16312), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1167)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_349_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8466_4_lut (.A(s_6_7), .B(n115), .C(n7_adj_476), .D(n7080), 
         .Z(n6_adj_935)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8466_4_lut.init = 16'h3022;
    LUT4 mux_308_i9_3_lut (.A(n18[8]), .B(instruction[8]), .C(n1339), 
         .Z(n1194[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i9_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_541_i12_3_lut_4_lut (.A(n22232), .B(n7908), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1168)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_541_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17472_2_lut (.A(instruction[15]), .B(instruction[14]), .Z(n20074)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17472_2_lut.init = 16'h6666;
    LUT4 i8561_4_lut (.A(n2340), .B(rst_n_in), .C(n2341), .D(n2323), 
         .Z(n1742[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8561_4_lut.init = 16'hc088;
    LUT4 PrioSelect_545_i12_3_lut_4_lut (.A(n22232), .B(n7908), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1169)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_545_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1818_3_lut_4_lut (.A(n22118), .B(n11714), .C(n7_adj_481), .D(n7_adj_500), 
         .Z(n10_adj_804)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1818_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1834_3_lut_4_lut (.A(n22118), .B(n11714), .C(n7_c), .D(n7_adj_479), 
         .Z(n10_adj_818)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1834_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_345_i13_3_lut_4_lut (.A(n22252), .B(n16312), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1170)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_345_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1850_3_lut_4_lut (.A(n22118), .B(n11714), .C(n7_adj_462), .D(n7_adj_481), 
         .Z(n10_adj_808)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1850_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_549_i12_3_lut_4_lut (.A(n22232), .B(n7908), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1171)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_549_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_308_i8_3_lut (.A(n18[7]), .B(instruction[7]), .C(n1339), 
         .Z(n1194[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i8_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_341_i13_3_lut_4_lut (.A(n22252), .B(n16312), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1172)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_341_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_337_i13_3_lut_4_lut (.A(n22252), .B(n16312), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1173)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_337_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1866_3_lut_4_lut (.A(n22118), .B(n11714), .C(n7_adj_609), .D(n7_c), 
         .Z(n10_adj_806)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1866_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_337_i14_3_lut_4_lut (.A(n22251), .B(n16312), .C(Z_N_387[1]), 
         .D(n13_adj_1173), .Z(n14_adj_977)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_337_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_525_i15_3_lut_4_lut (.A(n22232), .B(n7908), .C(n1108[0]), 
         .D(n5_adj_1174), .Z(n15_adj_985)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_525_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i8460_4_lut (.A(s_6_0), .B(n7), .C(n7_adj_2), .D(n7762), .Z(n2_adj_927)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8460_4_lut.init = 16'hceaa;
    LUT4 PrioSelect_553_i15_3_lut_4_lut (.A(n22232), .B(n7908), .C(n1108[7]), 
         .D(n9_adj_1175), .Z(n15_adj_1176)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_553_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_341_i14_3_lut_4_lut (.A(n22251), .B(n16312), .C(Z_N_387[2]), 
         .D(n13_adj_1172), .Z(n14_adj_993)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_341_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 instruction_17__I_0_532_i9_2_lut (.A(instruction[16]), .B(instruction[17]), 
         .Z(n9_adj_815)) /* synthesis lut_function=(A+!(B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(258[16:25])
    defparam instruction_17__I_0_532_i9_2_lut.init = 16'hbbbb;
    LUT4 PrioSelect_345_i14_3_lut_4_lut (.A(n22251), .B(n16312), .C(Z_N_387[3]), 
         .D(n13_adj_1170), .Z(n14_adj_989)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_345_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_adj_116 (.A(rst_n_in), .B(jp), .C(clk_in_c_enable_109), 
         .D(n14414), .Z(n1124)) /* synthesis lut_function=(A (B+!((D)+!C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_4_lut_adj_116.init = 16'h88a8;
    LUT4 i2_3_lut (.A(n20), .B(n11804), .C(instruction[17]), .Z(n14414)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 PrioSelect_349_i14_3_lut_4_lut (.A(n22251), .B(n16312), .C(Z_N_387[4]), 
         .D(n13_adj_1167), .Z(n14_adj_981)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_349_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_353_i14_3_lut_4_lut (.A(n22251), .B(n16312), .C(Z_N_387[5]), 
         .D(n13_adj_1166), .Z(n14_adj_990)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_353_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8560_4_lut (.A(n2338), .B(rst_n_in), .C(n2339), .D(n2323), 
         .Z(n1742[7])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8560_4_lut.init = 16'hc088;
    LUT4 i1882_3_lut_4_lut (.A(n22118), .B(n11714), .C(n7_adj_476), .D(n7_adj_462), 
         .Z(n10_adj_810)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1882_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_308_i7_3_lut (.A(n18[6]), .B(instruction[6]), .C(n1339), 
         .Z(n1194[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i7_3_lut.init = 16'hcaca;
    LUT4 i8559_4_lut (.A(n2336), .B(rst_n_in), .C(n2337), .D(n2323), 
         .Z(n1742[6])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8559_4_lut.init = 16'hc088;
    LUT4 i1898_3_lut_4_lut (.A(n22118), .B(n11714), .C(n7_adj_473), .D(n7_adj_609), 
         .Z(n10_adj_802)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1898_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3034_3_lut_4_lut (.A(n22233), .B(n7908), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1177)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i3034_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_357_i14_3_lut_4_lut (.A(n22251), .B(n16312), .C(Z_N_387[6]), 
         .D(n13_adj_1160), .Z(n14_adj_976)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_357_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_308_i6_3_lut (.A(n18[5]), .B(instruction[5]), .C(n1339), 
         .Z(n1194[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i6_3_lut.init = 16'hcaca;
    LUT4 i8451_4_lut (.A(s_5_0), .B(n10), .C(n10_adj_3), .D(n7762), 
         .Z(n2_adj_922)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8451_4_lut.init = 16'hceaa;
    LUT4 PrioSelect_333_i14_3_lut_4_lut (.A(n22251), .B(n16312), .C(Z_N_387[0]), 
         .D(n10_adj_1157), .Z(n14_adj_965)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_333_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_549_i13_3_lut_4_lut (.A(n22233), .B(n7908), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1178)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_549_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_361_i14_3_lut_4_lut (.A(n22251), .B(n16312), .C(Z_N_387[7]), 
         .D(n10_adj_1156), .Z(n14_adj_558)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_361_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_adj_117 (.A(instruction[14]), .B(instruction[12]), .Z(n4_adj_1039)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_117.init = 16'h4444;
    LUT4 i8558_4_lut (.A(n2334), .B(rst_n_in), .C(n2335), .D(n2323), 
         .Z(n1742[5])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8558_4_lut.init = 16'hc088;
    LUT4 mux_308_i5_3_lut (.A(n18[4]), .B(instruction[4]), .C(n1339), 
         .Z(n1194[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i5_3_lut.init = 16'hcaca;
    LUT4 i8557_4_lut (.A(n2332), .B(rst_n_in), .C(n2333), .D(n2323), 
         .Z(n1742[4])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8557_4_lut.init = 16'hc088;
    LUT4 PrioSelect_373_i11_3_lut_4_lut (.A(n22255), .B(n16312), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1179)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_373_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_308_i4_3_lut (.A(n18[3]), .B(instruction[3]), .C(n1339), 
         .Z(n1194[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i4_3_lut.init = 16'hcaca;
    LUT4 i8556_4_lut (.A(n2330), .B(rst_n_in), .C(n2331), .D(n2323), 
         .Z(n1742[3])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8556_4_lut.init = 16'hc088;
    LUT4 i8448_4_lut (.A(s_4_7), .B(n117), .C(n7_adj_476), .D(n7052), 
         .Z(n6_adj_914)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8448_4_lut.init = 16'h3022;
    PFUMX PrioSelect_109_i16 (.BLUT(n14_adj_1180), .ALUT(n15_adj_1181), 
          .C0(n16998), .Z(n16_adj_1182)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_237_i5_3_lut_4_lut (.A(n7762), .B(n22119), .C(n7_adj_479), 
         .D(n7_adj_473), .Z(n5_adj_1183)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_237_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i2042_3_lut_4_lut (.A(n7762), .B(n22119), .C(n7_adj_481), .D(n7_adj_500), 
         .Z(n10_adj_867)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2042_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_308_i3_3_lut (.A(n18[2]), .B(instruction[2]), .C(n1339), 
         .Z(n1194[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i3_3_lut.init = 16'hcaca;
    LUT4 i8555_4_lut (.A(n2328), .B(rst_n_in), .C(n2329), .D(n2323), 
         .Z(n1742[2])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8555_4_lut.init = 16'hc088;
    LUT4 mux_308_i2_3_lut (.A(n18[1]), .B(instruction[1]), .C(n1339), 
         .Z(n1194[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_308_i2_3_lut.init = 16'hcaca;
    LUT4 i8554_4_lut (.A(n2326), .B(rst_n_in), .C(n2327), .D(n2323), 
         .Z(n1742[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i8554_4_lut.init = 16'hc088;
    LUT4 i2058_3_lut_4_lut (.A(n7762), .B(n22119), .C(n7_c), .D(n7_adj_479), 
         .Z(n10_adj_874)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2058_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_545_i13_3_lut_4_lut (.A(n22233), .B(n7908), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1184)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_545_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_541_i13_3_lut_4_lut (.A(n22233), .B(n7908), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1185)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_541_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i8442_4_lut (.A(s_4_0), .B(n8), .C(n8_adj_4), .D(n7762), .Z(n2_adj_901)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8442_4_lut.init = 16'hceaa;
    LUT4 PrioSelect_369_i11_3_lut_4_lut (.A(n22255), .B(n16312), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1186)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_369_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i2074_3_lut_4_lut (.A(n7762), .B(n22119), .C(n7_adj_462), .D(n7_adj_481), 
         .Z(n10_adj_869)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2074_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_537_i13_3_lut_4_lut (.A(n22233), .B(n7908), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1187)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_537_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i8433_4_lut (.A(s_3_0), .B(n9), .C(n9_adj_1), .D(n11714), .Z(n2_adj_891)) /* synthesis lut_function=(A (B+((D)+!C))+!A !((D)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8433_4_lut.init = 16'haace;
    LUT4 PrioSelect_377_i11_3_lut_4_lut (.A(n22255), .B(n16312), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1188)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_377_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i6028_2_lut (.A(instruction[9]), .B(n8773), .Z(n8647)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i6028_2_lut.init = 16'h8888;
    LUT4 PrioSelect_381_i11_3_lut_4_lut (.A(n22255), .B(n16312), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1189)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_381_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_533_i13_3_lut_4_lut (.A(n22233), .B(n7908), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1190)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_533_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_385_i11_3_lut_4_lut (.A(n22255), .B(n16312), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1191)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_385_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_389_i11_3_lut_4_lut (.A(n22255), .B(n16312), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1192)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_389_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_529_i13_3_lut_4_lut (.A(n22233), .B(n7908), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1193)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_529_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i8430_4_lut (.A(s_2_7), .B(n16264), .C(n7_adj_476), .D(n16245), 
         .Z(n6_adj_884)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8430_4_lut.init = 16'h3022;
    LUT4 PrioSelect_393_i11_3_lut_4_lut (.A(n22253), .B(n16312), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1194)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_393_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i2090_3_lut_4_lut (.A(n7762), .B(n22119), .C(n7_adj_609), .D(n7_c), 
         .Z(n10_adj_868)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2090_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_365_i11_3_lut_4_lut (.A(n22253), .B(n16312), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1195)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_365_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i17522_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22258), .B(n16312), .C(n22255), 
         .D(n22253), .Z(n18306)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17522_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hccc8;
    LUT4 PrioSelect_365_i12_3_lut_4_lut (.A(n22258), .B(n16312), .C(Z_N_378[0]), 
         .D(n11_adj_1195), .Z(n12_adj_1196)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_365_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17593_2_lut_3_lut_4_lut (.A(n7908), .B(n22266), .C(n20194), 
         .D(n16392), .Z(n19361)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;
    defparam i17593_2_lut_3_lut_4_lut.init = 16'hf2f0;
    CCU2D add_21_13 (.A0(address[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pc[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14270), 
          .S0(n18[11]), .S1(n18[12]));   // f:/home/mini-mcu/step_fpga/mcu.v(217[27:35])
    defparam add_21_13.INIT0 = 16'h5aaa;
    defparam add_21_13.INIT1 = 16'h5aaa;
    defparam add_21_13.INJECT1_0 = "NO";
    defparam add_21_13.INJECT1_1 = "NO";
    LUT4 i17704_2_lut_3_lut_4_lut (.A(n7908), .B(n22266), .C(n20305), 
         .D(n11778), .Z(n18993)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;
    defparam i17704_2_lut_3_lut_4_lut.init = 16'hf0f2;
    LUT4 PrioSelect_393_i12_3_lut_4_lut (.A(n22258), .B(n16312), .C(Z_N_378[7]), 
         .D(n11_adj_1194), .Z(n12_adj_544)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_393_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_553_i10_3_lut_4_lut (.A(n22233), .B(n7908), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1197)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_553_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i8424_4_lut (.A(s_2_0), .B(n7), .C(n7_adj_2), .D(n11714), .Z(n2_adj_880)) /* synthesis lut_function=(A (B+((D)+!C))+!A !((D)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8424_4_lut.init = 16'haace;
    LUT4 PrioSelect_529_i14_3_lut_4_lut (.A(n22234), .B(n7908), .C(Z_N_387[1]), 
         .D(n13_adj_1193), .Z(n14_adj_1061)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_529_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_533_i14_3_lut_4_lut (.A(n22234), .B(n7908), .C(Z_N_387[2]), 
         .D(n13_adj_1190), .Z(n14_adj_1085)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_533_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_537_i14_3_lut_4_lut (.A(n22234), .B(n7908), .C(Z_N_387[3]), 
         .D(n13_adj_1187), .Z(n14_adj_1076)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_537_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_541_i14_3_lut_4_lut (.A(n22234), .B(n7908), .C(Z_N_387[4]), 
         .D(n13_adj_1185), .Z(n14_adj_1067)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_541_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 n2083_bdd_4_lut_17898 (.A(n22109), .B(n2085), .C(n7908), .D(n7726), 
         .Z(n21201)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam n2083_bdd_4_lut_17898.init = 16'h1fff;
    LUT4 PrioSelect_545_i14_3_lut_4_lut (.A(n22234), .B(n7908), .C(Z_N_387[5]), 
         .D(n13_adj_1184), .Z(n14_adj_1079)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_545_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17783_2_lut_3_lut_4_lut (.A(n22264), .B(n11778), .C(n20384), 
         .D(n7762), .Z(n17397)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17783_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i17527_2_lut_3_lut_4_lut (.A(n22264), .B(n11778), .C(n20128), 
         .D(n16312), .Z(n18282)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17527_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i8415_4_lut (.A(s_1_0), .B(n10), .C(n10_adj_3), .D(n11714), 
         .Z(n2_adj_855)) /* synthesis lut_function=(A (B+((D)+!C))+!A !((D)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8415_4_lut.init = 16'haace;
    LUT4 PrioSelect_141_i5_3_lut_4_lut (.A(n8647), .B(n11714), .C(n7_adj_479), 
         .D(n7_adj_473), .Z(n5_adj_1198)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_141_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2106_3_lut_4_lut (.A(n7762), .B(n22119), .C(n7_adj_476), .D(n7_adj_462), 
         .Z(n10_adj_873)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2106_3_lut_4_lut.init = 16'hf780;
    LUT4 i110_4_lut (.A(instruction[14]), .B(n1384), .C(instruction[16]), 
         .D(C_N_351[0]), .Z(n77)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i110_4_lut.init = 16'h3a30;
    LUT4 i17768_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n11778), .C(n7762), 
         .D(n22263), .Z(n17523)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+!(C)))) */ ;
    defparam i17768_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h1030;
    LUT4 i17753_2_lut_3_lut_4_lut (.A(n22264), .B(n11778), .C(n20354), 
         .D(n7762), .Z(n17546)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17753_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i17554_2_lut_3_lut_4_lut (.A(n22264), .B(n11778), .C(n20155), 
         .D(n16312), .Z(n18133)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17554_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 PrioSelect_549_i14_3_lut_4_lut (.A(n22234), .B(n7908), .C(Z_N_387[6]), 
         .D(n13_adj_1178), .Z(n14_adj_1058)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_549_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17691_2_lut_3_lut_4_lut (.A(n22264), .B(n11778), .C(n20292), 
         .D(n7908), .Z(n19018)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17691_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 PrioSelect_525_i14_3_lut_4_lut (.A(n22234), .B(n7908), .C(Z_N_387[0]), 
         .D(n10_adj_1177), .Z(n14_adj_984)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_525_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i2122_3_lut_4_lut (.A(n7762), .B(n22119), .C(n7_adj_473), .D(n7_adj_609), 
         .Z(n10_adj_866)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2122_3_lut_4_lut.init = 16'hf780;
    CCU2D add_632_7 (.A0(instruction[5]), .B0(n7_adj_609), .C0(instruction[11]), 
          .D0(n14_adj_705), .A1(instruction[6]), .B1(n7_adj_476), .C1(instruction[11]), 
          .D1(n14_adj_709), .CIN(n14263), .COUT(n14264), .S0(Z_N_367[5]), 
          .S1(Z_N_367[6]));   // f:/home/mini-mcu/step_fpga/mcu.v(263[59:70])
    defparam add_632_7.INIT0 = 16'h56a6;
    defparam add_632_7.INIT1 = 16'h56a6;
    defparam add_632_7.INJECT1_0 = "NO";
    defparam add_632_7.INJECT1_1 = "NO";
    LUT4 i17541_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n11778), .C(n16312), 
         .D(n22263), .Z(n18259)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+!(C)))) */ ;
    defparam i17541_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h1030;
    LUT4 PrioSelect_301_i5_3_lut_4_lut (.A(n7762), .B(n22118), .C(n7_adj_479), 
         .D(n7_adj_473), .Z(n5_adj_1091)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_301_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 Mux_7_i14_3_lut (.A(n19793), .B(n13_adj_739), .C(instruction[10]), 
         .Z(n14)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_7_i14_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_553_i14_3_lut_4_lut (.A(n22234), .B(n7908), .C(Z_N_387[7]), 
         .D(n10_adj_1197), .Z(n14_adj_1199)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_553_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17720_2_lut_3_lut_4_lut (.A(n22264), .B(n11778), .C(n20321), 
         .D(n7908), .Z(n18869)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17720_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 PrioSelect_369_i12_3_lut_4_lut (.A(n22254), .B(n16312), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1200)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_369_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17702_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n11778), .C(n7908), 
         .D(n22263), .Z(n18995)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+!(C)))) */ ;
    defparam i17702_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h1030;
    LUT4 PrioSelect_373_i12_3_lut_4_lut (.A(n22254), .B(n16312), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1201)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_373_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 Mux_6_i14_3_lut (.A(n19787), .B(n13_adj_516), .C(instruction[10]), 
         .Z(n14_adj_463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_6_i14_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_377_i12_3_lut_4_lut (.A(n22254), .B(n16312), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1202)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_377_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_381_i12_3_lut_4_lut (.A(n22254), .B(n16312), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1203)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_381_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i2298_3_lut_4_lut (.A(n7762), .B(n22118), .C(n7_adj_462), .D(n7_adj_481), 
         .Z(n10_adj_921)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2298_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_385_i12_3_lut_4_lut (.A(n22254), .B(n16312), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1204)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_385_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_389_i12_3_lut_4_lut (.A(n22254), .B(n16312), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1205)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_389_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_365_i15_3_lut_4_lut (.A(n22254), .B(n16312), .C(n1108[0]), 
         .D(n5_adj_1206), .Z(n15_adj_1083)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_365_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_393_i15_3_lut_4_lut (.A(n22254), .B(n16312), .C(n1108[7]), 
         .D(n9_adj_1010), .Z(n15_adj_540)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_393_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i2330_3_lut_4_lut (.A(n7762), .B(n22118), .C(n7_adj_476), .D(n7_adj_462), 
         .Z(n10_adj_930)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2330_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_393_i10_3_lut_4_lut (.A(n22259), .B(n16312), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1207)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_393_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i2474_3_lut_4_lut (.A(n22259), .B(n16312), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1208)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i2474_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_389_i13_3_lut_4_lut (.A(n22259), .B(n16312), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1209)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_389_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i8412_4_lut (.A(s_0_7), .B(n16265), .C(n7_adj_476), .D(n16253), 
         .Z(n6_adj_852)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8412_4_lut.init = 16'h3022;
    LUT4 PrioSelect_385_i13_3_lut_4_lut (.A(n22259), .B(n16312), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1210)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_385_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i17544_2_lut_rep_524_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n11778), 
         .C(n16312), .D(n22268), .Z(n22091)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+!(C)))) */ ;
    defparam i17544_2_lut_rep_524_3_lut_3_lut_4_lut_4_lut.init = 16'h1030;
    LUT4 PrioSelect_381_i13_3_lut_4_lut (.A(n22259), .B(n16312), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1211)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_381_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i2282_3_lut_4_lut (.A(n7762), .B(n22118), .C(n7_c), .D(n7_adj_479), 
         .Z(n10_adj_932)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2282_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_377_i13_3_lut_4_lut (.A(n22259), .B(n16312), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1212)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_377_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_373_i13_3_lut_4_lut (.A(n22259), .B(n16312), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1213)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_373_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_369_i13_3_lut_4_lut (.A(n22259), .B(n16312), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1214)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_369_i13_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_557_i16 (.BLUT(n14_adj_1215), .ALUT(n15_adj_1216), 
          .C0(n19574), .Z(n16_adj_1217)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17705_2_lut_rep_531_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n11778), 
         .C(n7908), .D(n22268), .Z(n22098)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+!(C)))) */ ;
    defparam i17705_2_lut_rep_531_3_lut_3_lut_4_lut_4_lut.init = 16'h1030;
    LUT4 and_168_i8_2_lut (.A(C_N_336[0]), .B(instruction[7]), .Z(Z_N_387[7])) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(351[112:121])
    defparam and_168_i8_2_lut.init = 16'h8888;
    LUT4 PrioSelect_369_i14_3_lut_4_lut (.A(n22257), .B(n16312), .C(Z_N_387[1]), 
         .D(n13_adj_1214), .Z(n14_adj_1002)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_369_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17771_2_lut_rep_520_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n11778), 
         .C(n7762), .D(n22268), .Z(n22087)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+!(C)))) */ ;
    defparam i17771_2_lut_rep_520_3_lut_3_lut_4_lut_4_lut.init = 16'h1030;
    LUT4 PrioSelect_373_i14_3_lut_4_lut (.A(n22257), .B(n16312), .C(Z_N_387[2]), 
         .D(n13_adj_1213), .Z(n14_adj_1006)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_373_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_377_i14_3_lut_4_lut (.A(n22257), .B(n16312), .C(Z_N_387[3]), 
         .D(n13_adj_1212), .Z(n14_adj_997)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_377_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_381_i14_3_lut_4_lut (.A(n22257), .B(n16312), .C(Z_N_387[4]), 
         .D(n13_adj_1211), .Z(n14_adj_1000)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_381_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 Mux_13_i15_3_lut (.A(n7_adj_473), .B(n14_adj_711), .C(instruction[11]), 
         .Z(C_N_336[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[71:78])
    defparam Mux_13_i15_3_lut.init = 16'hcaca;
    LUT4 i16465_3_lut (.A(n19633), .B(n19634), .C(instruction[7]), .Z(port_id_7__N_200[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16465_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_385_i14_3_lut_4_lut (.A(n22257), .B(n16312), .C(Z_N_387[5]), 
         .D(n13_adj_1210), .Z(n14_adj_1008)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_385_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_389_i14_3_lut_4_lut (.A(n22257), .B(n16312), .C(Z_N_387[6]), 
         .D(n13_adj_1209), .Z(n14_adj_1004)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_389_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_365_i14_3_lut_4_lut (.A(n22257), .B(n16312), .C(Z_N_387[0]), 
         .D(n10_adj_1208), .Z(n14_adj_1082)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_365_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i2314_3_lut_4_lut (.A(n7762), .B(n22118), .C(n7_adj_609), .D(n7_c), 
         .Z(n10_adj_913)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2314_3_lut_4_lut.init = 16'hf780;
    LUT4 i17701_2_lut_3_lut_4_lut (.A(n22264), .B(n7726), .C(n20302), 
         .D(n11714), .Z(n16994)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17701_2_lut_3_lut_4_lut.init = 16'hf0f4;
    LUT4 PrioSelect_393_i14_3_lut_4_lut (.A(n22257), .B(n16312), .C(Z_N_387[7]), 
         .D(n10_adj_1207), .Z(n14_adj_539)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_393_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17709_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n7726), .C(n7762), 
         .D(n22263), .Z(n17707)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17709_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i2346_3_lut_4_lut (.A(n7762), .B(n22118), .C(n7_adj_473), .D(n7_adj_609), 
         .Z(n10_adj_907)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2346_3_lut_4_lut.init = 16'hf780;
    LUT4 i17774_2_lut_3_lut_4_lut (.A(n22264), .B(n7726), .C(n20375), 
         .D(n11714), .Z(n16845)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17774_2_lut_3_lut_4_lut.init = 16'hf0f4;
    LUT4 i17696_2_lut_3_lut_4_lut (.A(n22264), .B(n7726), .C(n20297), 
         .D(n7762), .Z(n17730)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17696_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i17486_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n7726), .C(n16312), 
         .D(n22263), .Z(n18363)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17486_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i17745_2_lut_3_lut_4_lut (.A(n22264), .B(n7726), .C(n20346), 
         .D(n7762), .Z(n17581)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17745_2_lut_3_lut_4_lut.init = 16'hf4f0;
    CCU2D sub_131_add_2_9 (.A0(Z_N_378[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14281), .S0(n703[7]));   // f:/home/mini-mcu/step_fpga/mcu.v(281[61:73])
    defparam sub_131_add_2_9.INIT0 = 16'h5555;
    defparam sub_131_add_2_9.INIT1 = 16'h0000;
    defparam sub_131_add_2_9.INJECT1_0 = "NO";
    defparam sub_131_add_2_9.INJECT1_1 = "NO";
    LUT4 i17781_2_lut_3_lut_4_lut (.A(n22264), .B(n7726), .C(n20382), 
         .D(n16312), .Z(n18466)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17781_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i17665_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n7726), .C(n7908), 
         .D(n22263), .Z(n19179)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17665_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i2266_3_lut_4_lut (.A(n7762), .B(n22118), .C(n7_adj_481), .D(n7_adj_500), 
         .Z(n10_adj_911)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2266_3_lut_4_lut.init = 16'hf780;
    LUT4 i17494_2_lut_3_lut_4_lut (.A(n22264), .B(n7726), .C(n20095), 
         .D(n16312), .Z(n18317)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17494_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i17662_2_lut_3_lut_4_lut (.A(n22264), .B(n7726), .C(n20263), 
         .D(n7908), .Z(n19202)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17662_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i8406_4_lut (.A(s_0_0), .B(n8), .C(n8_adj_4), .D(n11714), .Z(n2)) /* synthesis lut_function=(A (B+((D)+!C))+!A !((D)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8406_4_lut.init = 16'haace;
    LUT4 i17714_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n7726), .C(n11714), 
         .D(n22263), .Z(n16971)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17714_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h040c;
    LUT4 PrioSelect_105_i11_3_lut_4_lut (.A(n22246), .B(n11714), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1218)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam PrioSelect_105_i11_3_lut_4_lut.init = 16'hfe10;
    LUT4 i17684_2_lut_3_lut_4_lut (.A(n22264), .B(n7726), .C(n20285), 
         .D(n7908), .Z(n19053)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17684_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 n2083_bdd_4_lut_17907 (.A(n22109), .B(n2085), .C(n7908), .D(n16392), 
         .Z(n21226)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam n2083_bdd_4_lut_17907.init = 16'h1fff;
    LUT4 PrioSelect_365_i5_3_lut_4_lut (.A(n22119), .B(n16312), .C(n14_adj_480), 
         .D(n14_adj_711), .Z(n5_adj_1206)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_365_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_77_i11_3_lut_4_lut (.A(n22246), .B(n11714), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1219)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam PrioSelect_77_i11_3_lut_4_lut.init = 16'hfe10;
    LUT4 PrioSelect_405_i11_3_lut_4_lut (.A(n22229), .B(n16312), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1220)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_405_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_401_i11_3_lut_4_lut (.A(n22229), .B(n16312), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1221)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_401_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_409_i11_3_lut_4_lut (.A(n22229), .B(n16312), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1222)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_409_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_413_i11_3_lut_4_lut (.A(n22229), .B(n16312), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1223)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_413_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_417_i11_3_lut_4_lut (.A(n22229), .B(n16312), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1224)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_417_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_421_i11_3_lut_4_lut (.A(n22229), .B(n16312), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1225)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_421_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i2490_3_lut_4_lut (.A(n22119), .B(n16312), .C(n14_adj_482), .D(n14_adj_501), 
         .Z(n10_adj_1003)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2490_3_lut_4_lut.init = 16'hf780;
    LUT4 i7_4_lut (.A(n16522), .B(Z_N_367[7]), .C(instruction[12]), .D(Z_N_367[0]), 
         .Z(n16_adj_848)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i7_4_lut.init = 16'h0010;
    LUT4 i13361_2_lut (.A(Z_N_367[5]), .B(Z_N_367[1]), .Z(n16522)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13361_2_lut.init = 16'heeee;
    LUT4 PrioSelect_425_i11_3_lut_4_lut (.A(n22230), .B(n16312), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1226)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_425_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_397_i11_3_lut_4_lut (.A(n22230), .B(n16312), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1227)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_397_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i13363_2_lut (.A(Z_N_367[4]), .B(Z_N_367[3]), .Z(n16524)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13363_2_lut.init = 16'heeee;
    LUT4 i2506_3_lut_4_lut (.A(n22119), .B(n16312), .C(n14), .D(n14_adj_480), 
         .Z(n10_adj_1007)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2506_3_lut_4_lut.init = 16'hf780;
    LUT4 i17762_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22231), .B(n16312), .C(n22229), 
         .D(n22230), .Z(n18642)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17762_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hccc8;
    LUT4 i2522_3_lut_4_lut (.A(n22119), .B(n16312), .C(n14_adj_463), .D(n14_adj_482), 
         .Z(n10_adj_998)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2522_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_497_i17_3_lut_4_lut (.A(n22266), .B(n16375), .C(in_port[1]), 
         .D(n16_adj_1228), .Z(n17)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_497_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1308_i3_4_lut_4_lut_then_4_lut (.A(st[0]), .B(st[1]), .C(n14459), 
         .D(st[2]), .Z(n22312)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[23:27])
    defparam mux_1308_i3_4_lut_4_lut_then_4_lut.init = 16'h7ffe;
    LUT4 PrioSelect_501_i17_3_lut_4_lut (.A(n22266), .B(n16375), .C(in_port[2]), 
         .D(n16_adj_1229), .Z(n17_adj_1230)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_501_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_425_i12_3_lut_4_lut (.A(n22231), .B(n16312), .C(Z_N_378[7]), 
         .D(n11_adj_1226), .Z(n12_adj_1231)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_425_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i13474_4_lut_4_lut_4_lut (.A(n22249), .B(n11714), .C(n22082), 
         .D(n8627), .Z(n16644)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B)) */ ;
    defparam i13474_4_lut_4_lut_4_lut.init = 16'hccce;
    LUT4 PrioSelect_397_i12_3_lut_4_lut (.A(n22231), .B(n16312), .C(Z_N_378[0]), 
         .D(n11_adj_1227), .Z(n12_adj_1232)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_397_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_505_i17_3_lut_4_lut (.A(n22266), .B(n16375), .C(in_port[3]), 
         .D(n16_adj_1233), .Z(n17_adj_1234)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_505_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i2538_3_lut_4_lut (.A(n22119), .B(n16312), .C(n14_adj_705), .D(n14), 
         .Z(n10_adj_1001)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2538_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_509_i17_3_lut_4_lut (.A(n22266), .B(n16375), .C(in_port[4]), 
         .D(n16_adj_1235), .Z(n17_adj_1236)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_509_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_513_i17_3_lut_4_lut (.A(n22266), .B(n16375), .C(in_port[5]), 
         .D(n16_adj_1237), .Z(n17_adj_1238)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_513_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8551_4_lut (.A(s_15_7), .B(n7934), .C(n13_adj_515), .D(n6928), 
         .Z(n6_adj_838)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8551_4_lut.init = 16'h3022;
    LUT4 i13622_4_lut_4_lut_4_lut (.A(n22249), .B(n11714), .C(n8_adj_5), 
         .D(n22101), .Z(n16792)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B)) */ ;
    defparam i13622_4_lut_4_lut_4_lut.init = 16'hccce;
    LUT4 PrioSelect_401_i12_3_lut_4_lut (.A(n22232), .B(n16312), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1240)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_401_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_517_i17_3_lut_4_lut (.A(n22266), .B(n16375), .C(in_port[6]), 
         .D(n16_adj_1241), .Z(n17_adj_1242)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_517_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i2554_3_lut_4_lut (.A(n22119), .B(n16312), .C(n14_adj_709), .D(n14_adj_463), 
         .Z(n10_adj_1009)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2554_3_lut_4_lut.init = 16'hf780;
    LUT4 i13381_2_lut (.A(instruction[8]), .B(instruction[9]), .Z(n11778)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13381_2_lut.init = 16'heeee;
    LUT4 PrioSelect_405_i12_3_lut_4_lut (.A(n22232), .B(n16312), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1243)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_405_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_409_i12_3_lut_4_lut (.A(n22232), .B(n16312), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1244)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_409_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_118 (.A(st_zc[1]), .B(n22283), .C(n22285), 
         .D(n22307), .Z(n1[2])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_118.init = 16'h0004;
    LUT4 PrioSelect_413_i12_3_lut_4_lut (.A(n22232), .B(n16312), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1245)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_413_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_417_i12_3_lut_4_lut (.A(n22232), .B(n16312), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1246)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_417_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i2570_3_lut_4_lut (.A(n22119), .B(n16312), .C(n14_adj_711), .D(n14_adj_705), 
         .Z(n10_adj_1005)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2570_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_421_i12_3_lut_4_lut (.A(n22232), .B(n16312), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1247)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_421_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 Mux_13_i14_3_lut (.A(n19754), .B(n13_adj_748), .C(instruction[10]), 
         .Z(n14_adj_711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[71:78])
    defparam Mux_13_i14_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_397_i15_3_lut_4_lut (.A(n22232), .B(n16312), .C(n1108[0]), 
         .D(n5_adj_713), .Z(n15_adj_961)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_397_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_429_i5_3_lut_4_lut (.A(n22118), .B(n16312), .C(n14_adj_480), 
         .D(n14_adj_711), .Z(n5_adj_1248)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_429_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_425_i15_3_lut_4_lut (.A(n22232), .B(n16312), .C(n1108[7]), 
         .D(n9_adj_1031), .Z(n15_adj_513)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_425_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i2762_3_lut_4_lut (.A(n22118), .B(n16312), .C(n14_adj_705), .D(n14), 
         .Z(n10_adj_1038)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2762_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_425_i10_3_lut_4_lut (.A(n22233), .B(n16312), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1249)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_425_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i2586_3_lut_4_lut (.A(n22233), .B(n16312), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1250)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i2586_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_421_i13_3_lut_4_lut (.A(n22233), .B(n16312), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1251)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_421_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i2778_3_lut_4_lut (.A(n22118), .B(n16312), .C(n14_adj_709), .D(n14_adj_463), 
         .Z(n10_adj_1046)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2778_3_lut_4_lut.init = 16'hf780;
    LUT4 i2714_3_lut_4_lut (.A(n22118), .B(n16312), .C(n14_adj_482), .D(n14_adj_501), 
         .Z(n10_adj_1035)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2714_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_417_i13_3_lut_4_lut (.A(n22233), .B(n16312), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1252)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_417_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 Mux_67_i14_3_lut (.A(n19796), .B(n5_adj_737), .C(instruction[10]), 
         .Z(n14_adj_501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(406[24:28])
    defparam Mux_67_i14_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_413_i13_3_lut_4_lut (.A(n22233), .B(n16312), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1253)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_413_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_409_i13_3_lut_4_lut (.A(n22233), .B(n16312), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1254)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_409_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i2730_3_lut_4_lut (.A(n22118), .B(n16312), .C(n14), .D(n14_adj_480), 
         .Z(n10_adj_1048)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2730_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_405_i13_3_lut_4_lut (.A(n22233), .B(n16312), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1255)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_405_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i2746_3_lut_4_lut (.A(n22118), .B(n16312), .C(n14_adj_463), .D(n14_adj_482), 
         .Z(n10_adj_1044)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2746_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_401_i13_3_lut_4_lut (.A(n22233), .B(n16312), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1256)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_401_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i17568_4_lut (.A(n22114), .B(n22116), .C(n22115), .D(n19532), 
         .Z(n20170)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17568_4_lut.init = 16'habaa;
    LUT4 PrioSelect_401_i14_3_lut_4_lut (.A(n22234), .B(n16312), .C(Z_N_387[1]), 
         .D(n13_adj_1256), .Z(n14_adj_1018)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_401_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17712_2_lut_rep_521_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n7726), 
         .C(n7762), .D(n22268), .Z(n22088)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17712_2_lut_rep_521_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 PrioSelect_405_i14_3_lut_4_lut (.A(n22234), .B(n16312), .C(Z_N_387[2]), 
         .D(n13_adj_1255), .Z(n14_adj_1030)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_405_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i2794_3_lut_4_lut (.A(n22118), .B(n16312), .C(n14_adj_711), .D(n14_adj_705), 
         .Z(n10_adj_1033)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2794_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_493_i5_3_lut_4_lut (.A(n22119), .B(n7908), .C(n13_adj_731), 
         .D(n14_adj_711), .Z(n5_adj_623)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_493_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i16342_4_lut (.A(n22108), .B(n22112), .C(n22113), .D(n213[15]), 
         .Z(n19532)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i16342_4_lut.init = 16'h5554;
    LUT4 i2938_3_lut_4_lut (.A(n22119), .B(n7908), .C(n13_adj_736), .D(n5_adj_737), 
         .Z(n10_adj_1257)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2938_3_lut_4_lut.init = 16'hf780;
    LUT4 i17480_2_lut_rep_525_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n7726), 
         .C(n16312), .D(n22268), .Z(n22092)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17480_2_lut_rep_525_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i17668_2_lut_rep_535_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n7726), 
         .C(n7908), .D(n22268), .Z(n22102)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17668_2_lut_rep_535_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i17717_2_lut_rep_517_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n7726), 
         .C(n11714), .D(n22268), .Z(n22084)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17717_2_lut_rep_517_3_lut_3_lut_4_lut_4_lut.init = 16'h040c;
    LUT4 i2954_3_lut_4_lut (.A(n22119), .B(n7908), .C(n13_adj_739), .D(n13_adj_731), 
         .Z(n10_adj_529)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2954_3_lut_4_lut.init = 16'hf780;
    LUT4 i8541_4_lut (.A(s_14_7), .B(n7933), .C(n13_adj_515), .D(n6914), 
         .Z(n6_adj_781)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8541_4_lut.init = 16'h3022;
    LUT4 PrioSelect_409_i14_3_lut_4_lut (.A(n22234), .B(n16312), .C(Z_N_387[3]), 
         .D(n13_adj_1254), .Z(n14_adj_1022)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_409_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i13413_3_lut_rep_654_4_lut (.A(n22270), .B(n22269), .C(n11916), 
         .D(n22271), .Z(n22221)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i13413_3_lut_rep_654_4_lut.init = 16'h8000;
    LUT4 i13390_2_lut_rep_694 (.A(n160), .B(n7646), .Z(n22261)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13390_2_lut_rep_694.init = 16'h8888;
    LUT4 i2970_3_lut_4_lut (.A(n22119), .B(n7908), .C(n13_adj_516), .D(n13_adj_736), 
         .Z(n10_c)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2970_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_413_i14_3_lut_4_lut (.A(n22234), .B(n16312), .C(Z_N_387[4]), 
         .D(n13_adj_1253), .Z(n14_adj_1021)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_413_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut_adj_119 (.A(n160), .B(n7646), .C(n22281), .D(instruction[3]), 
         .Z(n6928)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_119.init = 16'h0080;
    LUT4 PrioSelect_101_i13_3_lut_4_lut (.A(n22252), .B(n11714), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_661)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam PrioSelect_101_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 PrioSelect_417_i14_3_lut_4_lut (.A(n22234), .B(n16312), .C(Z_N_387[5]), 
         .D(n13_adj_1252), .Z(n14_adj_1027)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_417_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_120 (.A(st_zc[1]), .B(n22283), .C(n22282), 
         .D(n22307), .Z(n1[10])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(205[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_120.init = 16'h0040;
    LUT4 i1_2_lut_adj_121 (.A(n8789), .B(n8044), .Z(n6914)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_adj_121.init = 16'h8888;
    LUT4 PrioSelect_97_i13_3_lut_4_lut (.A(n22252), .B(n11714), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_659)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam PrioSelect_97_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 PrioSelect_105_i10_3_lut_4_lut (.A(n22252), .B(n11714), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_652)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam PrioSelect_105_i10_3_lut_4_lut.init = 16'hfe10;
    LUT4 PrioSelect_421_i14_3_lut_4_lut (.A(n22234), .B(n16312), .C(Z_N_387[6]), 
         .D(n13_adj_1251), .Z(n14_adj_1013)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_421_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_397_i14_3_lut_4_lut (.A(n22234), .B(n16312), .C(Z_N_387[0]), 
         .D(n10_adj_1250), .Z(n14_adj_960)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_397_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_425_i14_3_lut_4_lut (.A(n22234), .B(n16312), .C(Z_N_387[7]), 
         .D(n10_adj_1249), .Z(n14_adj_512)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_425_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i1466_3_lut_4_lut (.A(n22252), .B(n11714), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_648)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i1466_3_lut_4_lut.init = 16'hfe10;
    LUT4 PrioSelect_93_i13_3_lut_4_lut (.A(n22252), .B(n11714), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_655)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam PrioSelect_93_i13_3_lut_4_lut.init = 16'hfe10;
    CCU2D sub_131_add_2_7 (.A0(Z_N_378[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Z_N_378[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14280), .COUT(n14281), .S0(n703[5]), .S1(n703[6]));   // f:/home/mini-mcu/step_fpga/mcu.v(281[61:73])
    defparam sub_131_add_2_7.INIT0 = 16'h5555;
    defparam sub_131_add_2_7.INIT1 = 16'h5555;
    defparam sub_131_add_2_7.INJECT1_0 = "NO";
    defparam sub_131_add_2_7.INJECT1_1 = "NO";
    LUT4 i17646_4_lut_4_lut (.A(n22276), .B(n11778), .C(n11714), .D(n8050), 
         .Z(n9164)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i17646_4_lut_4_lut.init = 16'h0001;
    LUT4 PrioSelect_437_i11_3_lut_4_lut (.A(n22235), .B(n16312), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1258)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_437_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i17654_3_lut_rep_695 (.A(rst_n_in), .B(jp), .C(n4), .Z(clk_in_c_enable_159)) /* synthesis lut_function=(!(A (B+(C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i17654_3_lut_rep_695.init = 16'h5757;
    LUT4 i17460_2_lut_4_lut (.A(rst_n_in), .B(jp), .C(n4), .D(st_zc[0]), 
         .Z(n20062)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A !(D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i17460_2_lut_4_lut.init = 16'ha857;
    LUT4 PrioSelect_433_i11_3_lut_4_lut (.A(n22235), .B(n16312), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1259)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_433_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_89_i13_3_lut_4_lut (.A(n22252), .B(n11714), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_625)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam PrioSelect_89_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 i17592_4_lut (.A(n22120), .B(n22122), .C(n22121), .D(n19348), 
         .Z(n20194)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17592_4_lut.init = 16'habaa;
    LUT4 PrioSelect_85_i13_3_lut_4_lut (.A(n22252), .B(n11714), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_531)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam PrioSelect_85_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 PrioSelect_453_i11_3_lut_4_lut (.A(n22235), .B(n16312), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1260)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_453_i11_3_lut_4_lut.init = 16'hf780;
    CCU2D sub_131_add_2_5 (.A0(Z_N_378[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Z_N_378[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14279), .COUT(n14280), .S0(n703[3]), .S1(n703[4]));   // f:/home/mini-mcu/step_fpga/mcu.v(281[61:73])
    defparam sub_131_add_2_5.INIT0 = 16'h5555;
    defparam sub_131_add_2_5.INIT1 = 16'h5555;
    defparam sub_131_add_2_5.INJECT1_0 = "NO";
    defparam sub_131_add_2_5.INJECT1_1 = "NO";
    LUT4 i16158_4_lut (.A(n22107), .B(n22110), .C(n22111), .D(n213[14]), 
         .Z(n19348)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i16158_4_lut.init = 16'h5554;
    LUT4 PrioSelect_441_i11_3_lut_4_lut (.A(n22235), .B(n16312), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1261)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_441_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_81_i13_3_lut_4_lut (.A(n22252), .B(n11714), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_657)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam PrioSelect_81_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 i8532_4_lut (.A(s_13_7), .B(n7932), .C(n13_adj_515), .D(n6900), 
         .Z(n6_adj_721)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8532_4_lut.init = 16'h3022;
    LUT4 i2986_3_lut_4_lut (.A(n22119), .B(n7908), .C(n13_adj_744), .D(n13_adj_739), 
         .Z(n10_adj_1262)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2986_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_445_i11_3_lut_4_lut (.A(n22235), .B(n16312), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1263)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_445_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i5_4_lut (.A(instruction[16]), .B(n16558), .C(n22291), .D(n8_adj_830), 
         .Z(n7646)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i5_4_lut.init = 16'h2000;
    LUT4 PrioSelect_449_i11_3_lut_4_lut (.A(n22235), .B(n16312), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1264)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_449_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i13395_2_lut (.A(n16122), .B(instruction[15]), .Z(n16558)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13395_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_3_lut (.A(jp), .B(clk_in_c_enable_109), .C(rst_n_in), 
         .Z(n16409)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 st_1__bdd_4_lut (.A(st[1]), .B(st[2]), .C(n14459), .D(st[0]), 
         .Z(n21644)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (C+(D))+!B !(C+(D))))) */ ;
    defparam st_1__bdd_4_lut.init = 16'h6cc9;
    LUT4 i601_2_lut_rep_723_2_lut (.A(jp), .B(rst_n_in), .Z(clk_in_c_enable_115)) /* synthesis lut_function=(!(A+!(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i601_2_lut_rep_723_2_lut.init = 16'h4444;
    LUT4 PrioSelect_457_i11_3_lut_4_lut (.A(n22236), .B(n16312), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1265)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_457_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_429_i11_3_lut_4_lut (.A(n22236), .B(n16312), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1266)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_429_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i8186_2_lut_rep_733 (.A(rst_n_in), .B(jp), .Z(n22300)) /* synthesis lut_function=(A (B)) */ ;
    defparam i8186_2_lut_rep_733.init = 16'h8888;
    LUT4 mux_1308_i3_4_lut_4_lut_else_4_lut (.A(st[0]), .B(st[1]), .C(n14459), 
         .D(st[2]), .Z(n22311)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[23:27])
    defparam mux_1308_i3_4_lut_4_lut_else_4_lut.init = 16'h8001;
    LUT4 i17524_2_lut_2_lut_3_lut (.A(rst_n_in), .B(jp), .C(clk_in_c_enable_109), 
         .Z(clk_in_c_enable_173)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i17524_2_lut_2_lut_3_lut.init = 16'h7070;
    LUT4 rst_n_I_0_1_lut_rep_734 (.A(rst_n_in), .Z(n22301)) /* synthesis lut_function=(!(A)) */ ;   // f:/home/mini-mcu/step_fpga/divide.v(34[7:13])
    defparam rst_n_I_0_1_lut_rep_734.init = 16'h5555;
    LUT4 i17725_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22237), .B(n16312), .C(n22235), 
         .D(n22236), .Z(n18826)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17725_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hccc8;
    LUT4 i1372_2_lut_2_lut (.A(rst_n_in), .B(jp), .Z(n2730)) /* synthesis lut_function=((B)+!A) */ ;   // f:/home/mini-mcu/step_fpga/divide.v(34[7:13])
    defparam i1372_2_lut_2_lut.init = 16'hdddd;
    LUT4 PrioSelect_429_i12_3_lut_4_lut (.A(n22237), .B(n16312), .C(Z_N_378[0]), 
         .D(n11_adj_1266), .Z(n12_adj_1267)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_429_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i13415_4_lut (.A(instruction[4]), .B(instruction[6]), .C(instruction[5]), 
         .D(instruction[7]), .Z(n16122)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13415_4_lut.init = 16'hfffe;
    LUT4 PrioSelect_457_i12_3_lut_4_lut (.A(n22237), .B(n16312), .C(Z_N_378[7]), 
         .D(n11_adj_1265), .Z(n12)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_457_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i159_4_lut_4_lut (.A(rst_n_in), .B(\cnt_p[22] ), .C(\cnt_p[23] ), 
         .D(n14409), .Z(n857)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;   // f:/home/mini-mcu/step_fpga/divide.v(34[7:13])
    defparam i159_4_lut_4_lut.init = 16'hf5d5;
    LUT4 mux_1307_i2_4_lut_4_lut_4_lut (.A(st_zc[2]), .B(st_zc[1]), .C(st_zc[0]), 
         .D(clk_in_c_enable_109), .Z(n2634[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(206[26:38])
    defparam mux_1307_i2_4_lut_4_lut_4_lut.init = 16'ha96a;
    LUT4 i3002_3_lut_4_lut (.A(n22119), .B(n7908), .C(n13_adj_515), .D(n13_adj_516), 
         .Z(n10_adj_1268)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i3002_3_lut_4_lut.init = 16'hf780;
    LUT4 i3018_3_lut_4_lut (.A(n22119), .B(n7908), .C(n13_adj_748), .D(n13_adj_744), 
         .Z(n10_adj_1269)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i3018_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_516 (.A(n8773), .B(n8044), .Z(n22083)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1_2_lut_rep_516.init = 16'h8888;
    LUT4 PrioSelect_525_i5_3_lut_4_lut (.A(n8773), .B(n8044), .C(n13_adj_731), 
         .D(n14_adj_711), .Z(n5_adj_1174)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_525_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_717_3_lut_3_lut_4_lut (.A(rst_n_in), .B(jp), .C(st_zc[0]), 
         .D(clk_in_c_enable_109), .Z(n22284)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_2_lut_rep_717_3_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 n2083_bdd_4_lut_17922 (.A(n22109), .B(n2085), .C(n7908), .D(n7876), 
         .Z(n21255)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam n2083_bdd_4_lut_17922.init = 16'h1fff;
    LUT4 i1_2_lut_rep_716_3_lut_3_lut_4_lut (.A(rst_n_in), .B(jp), .C(st_zc[0]), 
         .D(clk_in_c_enable_109), .Z(n22283)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_2_lut_rep_716_3_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i17689_4_lut (.A(n22211), .B(n22213), .C(n22212), .D(n213[12]), 
         .Z(n19022)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17689_4_lut.init = 16'haaab;
    LUT4 i3050_3_lut_4_lut (.A(n8773), .B(n8044), .C(n13_adj_736), .D(n5_adj_737), 
         .Z(n10_adj_1062)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i3050_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_724_3_lut (.A(rst_n_in), .B(jp), .C(clk_in_c_enable_109), 
         .Z(n22291)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_2_lut_rep_724_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_122 (.A(rst_n_in), .B(jp), .C(n6978), 
         .D(clk_in_c_enable_109), .Z(creg_N_407)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_2_lut_3_lut_4_lut_adj_122.init = 16'h0200;
    LUT4 i8844_2_lut_rep_701_3_lut_3_lut_4_lut (.A(clk_in_c_enable_174), .B(instruction[15]), 
         .C(n9_adj_707), .D(n8_adj_708), .Z(n22268)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i8844_2_lut_rep_701_3_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i3066_3_lut_4_lut (.A(n8773), .B(n8044), .C(n13_adj_739), .D(n13_adj_731), 
         .Z(n10_adj_1086)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i3066_3_lut_4_lut.init = 16'hf780;
    LUT4 i1706_3_lut_4_lut (.A(n8647), .B(n11714), .C(n7_adj_481), .D(n7_adj_500), 
         .Z(n10_adj_784)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1706_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3082_3_lut_4_lut (.A(n8773), .B(n8044), .C(n13_adj_516), .D(n13_adj_736), 
         .Z(n10_adj_1077)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i3082_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_553_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n7908), 
         .D(n16392), .Z(n22120)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_553_3_lut_4_lut.init = 16'h1000;
    LUT4 i17520_4_lut_rep_736 (.A(enable_intr_flag), .B(intr_f[0]), .C(intr_f[2]), 
         .D(intr_f[1]), .Z(clk_in_c_enable_109)) /* synthesis lut_function=((B (C (D))+!B (C+!(D)))+!A) */ ;
    defparam i17520_4_lut_rep_736.init = 16'hf577;
    LUT4 i3098_3_lut_4_lut (.A(n8773), .B(n8044), .C(n13_adj_744), .D(n13_adj_739), 
         .Z(n10_adj_1068)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i3098_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_572_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n11714), 
         .D(n16392), .Z(n22139)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_572_3_lut_4_lut.init = 16'h0100;
    LUT4 i1722_3_lut_4_lut (.A(n8647), .B(n11714), .C(n7_c), .D(n7_adj_479), 
         .Z(n10_adj_798)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1722_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_596_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n7762), 
         .D(n16392), .Z(n22163)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_596_3_lut_4_lut.init = 16'h1000;
    LUT4 i1074_2_lut_rep_737 (.A(st_zc[1]), .B(st_zc[0]), .Z(n22304)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(206[26:38])
    defparam i1074_2_lut_rep_737.init = 16'h6666;
    LUT4 i1_2_lut_rep_620_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n16312), 
         .D(n16392), .Z(n22187)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_620_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_547_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n7908), 
         .D(n7876), .Z(n22114)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_547_3_lut_4_lut.init = 16'h1000;
    LUT4 i3114_3_lut_4_lut (.A(n8773), .B(n8044), .C(n13_adj_515), .D(n13_adj_516), 
         .Z(n10_adj_1080)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i3114_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_578_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n11714), 
         .D(n7876), .Z(n22145)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_578_3_lut_4_lut.init = 16'h0100;
    LUT4 i3130_3_lut_4_lut (.A(n8773), .B(n8044), .C(n13_adj_748), .D(n13_adj_744), 
         .Z(n10_adj_1059)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i3130_3_lut_4_lut.init = 16'hf780;
    LUT4 i13502_4_lut_4_lut (.A(n22123), .B(n22126), .C(n22124), .D(n22125), 
         .Z(n16672)) /* synthesis lut_function=(!(A (D)+!A (B (C+(D))+!B (D)))) */ ;
    defparam i13502_4_lut_4_lut.init = 16'h00bf;
    LUT4 i17550_4_lut_4_lut (.A(n22129), .B(n16672), .C(n22128), .D(n22127), 
         .Z(n20152)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B (D))) */ ;
    defparam i17550_4_lut_4_lut.init = 16'hff40;
    LUT4 PrioSelect_81_i17_3_lut (.A(n16_adj_1270), .B(in_port[1]), .C(n9164), 
         .Z(n17_adj_944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_81_i17_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_602_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n7762), 
         .D(n7876), .Z(n22169)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_602_3_lut_4_lut.init = 16'h1000;
    LUT4 i17483_4_lut_4_lut (.A(n22129), .B(n22126), .C(n22128), .D(n22127), 
         .Z(n16814)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B (D))) */ ;
    defparam i17483_4_lut_4_lut.init = 16'hff40;
    LUT4 i1_2_lut_rep_626_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n16312), 
         .D(n7876), .Z(n22193)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_626_3_lut_4_lut.init = 16'h1000;
    LUT4 PrioSelect_85_i17_3_lut (.A(n16_adj_1271), .B(in_port[2]), .C(n9164), 
         .Z(n17_adj_934)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_85_i17_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_608_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n16312), 
         .D(n11778), .Z(n22175)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_608_3_lut_4_lut.init = 16'h0010;
    CCU2D sub_131_add_2_3 (.A0(Z_N_378[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Z_N_378[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14278), .COUT(n14279), .S0(n703[1]), .S1(n703[2]));   // f:/home/mini-mcu/step_fpga/mcu.v(281[61:73])
    defparam sub_131_add_2_3.INIT0 = 16'h5555;
    defparam sub_131_add_2_3.INIT1 = 16'h5555;
    defparam sub_131_add_2_3.INJECT1_0 = "NO";
    defparam sub_131_add_2_3.INJECT1_1 = "NO";
    LUT4 PrioSelect_89_i17_3_lut (.A(n16_adj_1272), .B(in_port[3]), .C(n9164), 
         .Z(n17_adj_925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_89_i17_3_lut.init = 16'hcaca;
    LUT4 i1120_2_lut_rep_738 (.A(st[1]), .B(st[0]), .Z(n22305)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(284[52:61])
    defparam i1120_2_lut_rep_738.init = 16'h8888;
    LUT4 i1045_2_lut_3_lut (.A(st[1]), .B(st[0]), .C(st[2]), .Z(stack_N_397[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(284[52:61])
    defparam i1045_2_lut_3_lut.init = 16'h7878;
    LUT4 PrioSelect_93_i17_3_lut (.A(n16_adj_1273), .B(in_port[4]), .C(n9164), 
         .Z(n17_adj_917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_93_i17_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_584_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n7762), 
         .D(n11778), .Z(n22151)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_584_3_lut_4_lut.init = 16'h0010;
    LUT4 PrioSelect_97_i17_3_lut (.A(n16_adj_1274), .B(in_port[5]), .C(n9164), 
         .Z(n17_adj_904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_97_i17_3_lut.init = 16'hcaca;
    LUT4 i1052_2_lut_rep_721_3_lut_4_lut (.A(st[1]), .B(st[0]), .C(st[3]), 
         .D(st[2]), .Z(n22288)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(284[52:61])
    defparam i1052_2_lut_rep_721_3_lut_4_lut.init = 16'h78f0;
    LUT4 Mux_67_i15_3_lut (.A(n7_adj_500), .B(n14_adj_501), .C(instruction[11]), 
         .Z(out_port_7__N_217[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(406[24:28])
    defparam Mux_67_i15_3_lut.init = 16'hcaca;
    LUT4 Mux_9_i15_3_lut (.A(n7_adj_479), .B(n14_adj_480), .C(instruction[11]), 
         .Z(s_N_294[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_9_i15_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_101_i17_3_lut (.A(n16_adj_1275), .B(in_port[6]), .C(n9164), 
         .Z(n17_adj_890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_101_i17_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_644_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n7908), 
         .D(n11778), .Z(n22211)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_644_3_lut_4_lut.init = 16'h0010;
    LUT4 Mux_8_i15_3_lut (.A(n7_adj_481), .B(n14_adj_482), .C(instruction[11]), 
         .Z(s_N_294[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_8_i15_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_566_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n11714), 
         .D(n7726), .Z(n22133)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_566_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_590_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n7762), 
         .D(n7726), .Z(n22157)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_590_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_614_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n16312), 
         .D(n7726), .Z(n22181)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_614_3_lut_4_lut.init = 16'h1000;
    LUT4 Mux_7_i15_3_lut (.A(n7_c), .B(n14), .C(instruction[11]), .Z(s_N_294[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_7_i15_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_647_3_lut_4_lut (.A(n10_adj_698), .B(n22277), .C(n7908), 
         .D(n7726), .Z(n22214)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_647_3_lut_4_lut.init = 16'h1000;
    LUT4 PrioSelect_117_i11_3_lut_4_lut (.A(n22255), .B(n11714), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1276)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_117_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1188_2_lut_rep_739 (.A(st_zc[1]), .B(st_zc[0]), .Z(n22306)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(376[120:132])
    defparam i1188_2_lut_rep_739.init = 16'h8888;
    LUT4 PrioSelect_445_i12_3_lut_4_lut (.A(n22238), .B(n16312), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1277)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_445_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_113_i11_3_lut_4_lut (.A(n22255), .B(n11714), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1278)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_113_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 Mux_8_i14_3_lut (.A(n19742), .B(n13_adj_736), .C(instruction[10]), 
         .Z(n14_adj_482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_8_i14_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_449_i12_3_lut_4_lut (.A(n22238), .B(n16312), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1279)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_449_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1081_2_lut_rep_740 (.A(st_zc[1]), .B(st_zc[0]), .C(st_zc[2]), 
         .Z(n22307)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(376[120:132])
    defparam i1081_2_lut_rep_740.init = 16'h7878;
    LUT4 PrioSelect_433_i12_3_lut_4_lut (.A(n22238), .B(n16312), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1280)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_433_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_437_i12_3_lut_4_lut (.A(n22238), .B(n16312), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1281)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_437_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 Mux_9_i14_3_lut (.A(n19748), .B(n13_adj_731), .C(instruction[10]), 
         .Z(n14_adj_480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_9_i14_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_121_i11_3_lut_4_lut (.A(n22255), .B(n11714), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1282)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_121_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_adj_123 (.A(instruction[13]), .B(instruction[14]), .Z(n48)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_2_lut_adj_123.init = 16'h8888;
    LUT4 PrioSelect_441_i12_3_lut_4_lut (.A(n22238), .B(n16312), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1283)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_441_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_453_i12_3_lut_4_lut (.A(n22238), .B(n16312), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1284)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_453_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_429_i15_3_lut_4_lut (.A(n22238), .B(n16312), .C(n1108[0]), 
         .D(n5_adj_1248), .Z(n15_adj_1025)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_429_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_125_i11_3_lut_4_lut (.A(n22255), .B(n11714), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1285)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_125_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_457_i15_3_lut_4_lut (.A(n22238), .B(n16312), .C(n1108[7]), 
         .D(n9_adj_1050), .Z(n15_adj_492)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_457_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_129_i11_3_lut_4_lut (.A(n22255), .B(n11714), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1286)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_129_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_457_i10_3_lut_4_lut (.A(n22239), .B(n16312), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1287)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_457_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i2698_3_lut_4_lut (.A(n22239), .B(n16312), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1288)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i2698_3_lut_4_lut.init = 16'hf780;
    LUT4 i1139_2_lut_3_lut_4_lut (.A(st[1]), .B(st[0]), .C(st[3]), .D(st[2]), 
         .Z(n8_adj_1289)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(284[52:61])
    defparam i1139_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 PrioSelect_453_i13_3_lut_4_lut (.A(n22239), .B(n16312), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1290)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_453_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_449_i13_3_lut_4_lut (.A(n22239), .B(n16312), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1291)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_449_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_445_i13_3_lut_4_lut (.A(n22239), .B(n16312), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1292)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_445_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_441_i13_3_lut_4_lut (.A(n22239), .B(n16312), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1293)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_441_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_437_i13_3_lut_4_lut (.A(n22239), .B(n16312), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1294)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_437_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_433_i13_3_lut_4_lut (.A(n22239), .B(n16312), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1295)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_433_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_445_i14_3_lut_4_lut (.A(n22240), .B(n16312), .C(Z_N_387[4]), 
         .D(n13_adj_1292), .Z(n14_adj_1037)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_445_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_133_i11_3_lut_4_lut (.A(n22255), .B(n11714), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1296)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_133_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_449_i14_3_lut_4_lut (.A(n22240), .B(n16312), .C(Z_N_387[5]), 
         .D(n13_adj_1291), .Z(n14_adj_1045)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_449_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_433_i14_3_lut_4_lut (.A(n22240), .B(n16312), .C(Z_N_387[1]), 
         .D(n13_adj_1295), .Z(n14_adj_1034)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_433_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_437_i14_3_lut_4_lut (.A(n22240), .B(n16312), .C(Z_N_387[2]), 
         .D(n13_adj_1294), .Z(n14_adj_1047)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_437_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_441_i14_3_lut_4_lut (.A(n22240), .B(n16312), .C(Z_N_387[3]), 
         .D(n13_adj_1293), .Z(n14_adj_1043)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_441_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_453_i14_3_lut_4_lut (.A(n22240), .B(n16312), .C(Z_N_387[6]), 
         .D(n13_adj_1290), .Z(n14_adj_1032)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_453_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_429_i14_3_lut_4_lut (.A(n22240), .B(n16312), .C(Z_N_387[0]), 
         .D(n10_adj_1288), .Z(n14_adj_1024)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_429_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_457_i14_3_lut_4_lut (.A(n22240), .B(n16312), .C(Z_N_387[7]), 
         .D(n10_adj_1287), .Z(n14_adj_491)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_457_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_536_3_lut_4_lut (.A(n8050), .B(n22276), .C(n7876), 
         .D(n11714), .Z(n22103)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_536_3_lut_4_lut.init = 16'h0010;
    LUT4 PrioSelect_529_i17_3_lut_4_lut (.A(n16392), .B(n22247), .C(in_port[1]), 
         .D(n16_adj_1297), .Z(n17_adj_1298)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_529_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_533_i17_3_lut_4_lut (.A(n16392), .B(n22247), .C(in_port[2]), 
         .D(n16_adj_1299), .Z(n17_adj_1300)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_533_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_537_i17_3_lut_4_lut (.A(n16392), .B(n22247), .C(in_port[3]), 
         .D(n16_adj_1301), .Z(n17_adj_1302)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_537_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_537_3_lut_4_lut (.A(n8050), .B(n22276), .C(n16392), 
         .D(n11714), .Z(n22104)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_537_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_538_3_lut_4_lut (.A(n8050), .B(n22276), .C(n7726), 
         .D(n11714), .Z(n22105)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_538_3_lut_4_lut.init = 16'h0010;
    LUT4 PrioSelect_137_i11_3_lut_4_lut (.A(n22253), .B(n11714), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1303)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_137_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_109_i11_3_lut_4_lut (.A(n22253), .B(n11714), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1304)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_109_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17569_2_lut_3_lut_4_lut (.A(n8050), .B(n22276), .C(n20170), 
         .D(n22281), .Z(n19545)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17569_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 PrioSelect_541_i17_3_lut_4_lut (.A(n16392), .B(n22247), .C(in_port[4]), 
         .D(n16_adj_1305), .Z(n17_adj_1306)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_541_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_545_i17_3_lut_4_lut (.A(n16392), .B(n22247), .C(in_port[5]), 
         .D(n16_adj_1307), .Z(n17_adj_1308)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_545_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_630_3_lut_4_lut (.A(n8050), .B(n22276), .C(n7876), 
         .D(n16312), .Z(n22197)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_630_3_lut_4_lut.init = 16'h1000;
    LUT4 PrioSelect_549_i17_3_lut_4_lut (.A(n16392), .B(n22247), .C(in_port[6]), 
         .D(n16_adj_1309), .Z(n17_adj_1310)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_549_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_632_3_lut_4_lut (.A(n8050), .B(n22276), .C(n16392), 
         .D(n16312), .Z(n22199)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_632_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_633_3_lut_4_lut (.A(n8050), .B(n22276), .C(n7726), 
         .D(n16312), .Z(n22200)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_633_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_634_3_lut_4_lut (.A(n8050), .B(n22276), .C(n11778), 
         .D(n16312), .Z(n22201)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_634_3_lut_4_lut.init = 16'h0100;
    LUT4 PrioSelect_433_i17_3_lut_4_lut (.A(n7876), .B(n22242), .C(in_port[1]), 
         .D(n16_adj_1311), .Z(n17_adj_511)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_433_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_635_3_lut_4_lut (.A(n8050), .B(n22276), .C(n7876), 
         .D(n7762), .Z(n22202)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_635_3_lut_4_lut.init = 16'h1000;
    LUT4 PrioSelect_437_i17_3_lut_4_lut (.A(n7876), .B(n22242), .C(in_port[2]), 
         .D(n16_adj_1312), .Z(n17_adj_509)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_437_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_441_i17_3_lut_4_lut (.A(n7876), .B(n22242), .C(in_port[3]), 
         .D(n16_adj_1313), .Z(n17_adj_507)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_441_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_445_i17_3_lut_4_lut (.A(n7876), .B(n22242), .C(in_port[4]), 
         .D(n16_adj_1314), .Z(n17_adj_505)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_445_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_449_i17_3_lut_4_lut (.A(n7876), .B(n22242), .C(in_port[5]), 
         .D(n16_adj_1315), .Z(n17_adj_503)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_449_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_453_i17_3_lut_4_lut (.A(n7876), .B(n22242), .C(in_port[6]), 
         .D(n16_adj_1316), .Z(n17_adj_499)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_453_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut_adj_124 (.A(n22221), .B(n22280), .C(n15_adj_833), 
         .D(n7908), .Z(clk_in_c_enable_100)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_124.init = 16'hf400;
    LUT4 i17708_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22258), .B(n11714), .C(n22255), 
         .D(n22253), .Z(n16986)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17708_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3332;
    LUT4 i1_2_lut_rep_636_3_lut_4_lut (.A(n8050), .B(n22276), .C(n16392), 
         .D(n7762), .Z(n22203)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_636_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_637_3_lut_4_lut (.A(n8050), .B(n22276), .C(n7726), 
         .D(n7762), .Z(n22204)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_637_3_lut_4_lut.init = 16'h1000;
    LUT4 PrioSelect_109_i12_3_lut_4_lut (.A(n22258), .B(n11714), .C(Z_N_378[0]), 
         .D(n11_adj_1304), .Z(n12_adj_1317)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_109_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_137_i12_3_lut_4_lut (.A(n22258), .B(n11714), .C(Z_N_378[7]), 
         .D(n11_adj_1303), .Z(n12_adj_846)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_137_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_401_i17_3_lut_4_lut (.A(n16392), .B(n22242), .C(in_port[1]), 
         .D(n16_adj_1318), .Z(n17_adj_538)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_401_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_405_i17_3_lut_4_lut (.A(n16392), .B(n22242), .C(in_port[2]), 
         .D(n16_adj_1319), .Z(n17_adj_536)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_405_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_409_i17_3_lut_4_lut (.A(n16392), .B(n22242), .C(in_port[3]), 
         .D(n16_adj_1320), .Z(n17_adj_534)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_409_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_413_i17_3_lut_4_lut (.A(n16392), .B(n22242), .C(in_port[4]), 
         .D(n16_adj_1321), .Z(n17_adj_526)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_413_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1286_1_lut (.A(instruction[14]), .Z(n13_adj_844)) /* synthesis lut_function=(!(A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(216[16:21])
    defparam i1286_1_lut.init = 16'h5555;
    LUT4 i1285_1_lut (.A(instruction[16]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(216[16:21])
    defparam i1285_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_639_3_lut_4_lut (.A(n8050), .B(n22276), .C(n11778), 
         .D(n7762), .Z(n22206)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_639_3_lut_4_lut.init = 16'h0100;
    LUT4 PrioSelect_417_i17_3_lut_4_lut (.A(n16392), .B(n22242), .C(in_port[5]), 
         .D(n16_adj_1322), .Z(n17_adj_524)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_417_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i17642_4_lut_4_lut (.A(n22129), .B(n16652), .C(n22128), .D(n22127), 
         .Z(n16662)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i17642_4_lut_4_lut.init = 16'hffef;
    LUT4 i13630_4_lut_4_lut (.A(n22123), .B(n16792), .C(n22124), .D(n22125), 
         .Z(n16800)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i13630_4_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_629_3_lut_4_lut (.A(n8050), .B(n22276), .C(n16392), 
         .D(n7908), .Z(n22196)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_629_3_lut_4_lut.init = 16'h1000;
    LUT4 PrioSelect_421_i17_3_lut_4_lut (.A(n16392), .B(n22242), .C(in_port[6]), 
         .D(n16_adj_1323), .Z(n17_adj_522)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_421_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_369_i17_3_lut_4_lut (.A(n7726), .B(n22242), .C(in_port[1]), 
         .D(n16_adj_1324), .Z(n17_adj_557)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_369_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_373_i17_3_lut_4_lut (.A(n7726), .B(n22242), .C(in_port[2]), 
         .D(n16_adj_1325), .Z(n17_adj_555)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_373_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_377_i17_3_lut_4_lut (.A(n7726), .B(n22242), .C(in_port[3]), 
         .D(n16_adj_1326), .Z(n17_adj_553)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_377_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_381_i17_3_lut_4_lut (.A(n7726), .B(n22242), .C(in_port[4]), 
         .D(n16_adj_1327), .Z(n17_adj_551)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_381_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_385_i17_3_lut_4_lut (.A(n7726), .B(n22242), .C(in_port[5]), 
         .D(n16_adj_1328), .Z(n17_adj_549)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_385_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_389_i17_3_lut_4_lut (.A(n7726), .B(n22242), .C(in_port[6]), 
         .D(n16_adj_1329), .Z(n17_adj_547)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_389_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_642_3_lut_4_lut (.A(n8050), .B(n22276), .C(n11778), 
         .D(n7908), .Z(n22209)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_642_3_lut_4_lut.init = 16'h0100;
    LUT4 PrioSelect_113_i12_3_lut_4_lut (.A(n22254), .B(n11714), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1330)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_113_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17667_2_lut_3_lut_4_lut (.A(n8050), .B(n22276), .C(n20268), 
         .D(n16375), .Z(n19177)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17667_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i1_2_lut_rep_555_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n7908), 
         .D(n16392), .Z(n22122)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_555_3_lut_4_lut.init = 16'h1000;
    LUT4 i17703_4_lut (.A(n22211), .B(n22213), .C(n22212), .D(n18980), 
         .Z(n20305)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17703_4_lut.init = 16'habaa;
    LUT4 i15790_4_lut (.A(n22210), .B(n22208), .C(n22207), .D(n213[12]), 
         .Z(n18980)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15790_4_lut.init = 16'h5554;
    LUT4 PrioSelect_337_i17_3_lut_4_lut (.A(n11778), .B(n22242), .C(in_port[1]), 
         .D(n16_adj_1331), .Z(n17_adj_573)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_337_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_341_i17_3_lut_4_lut (.A(n11778), .B(n22242), .C(in_port[2]), 
         .D(n16_adj_1332), .Z(n17_adj_571)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_341_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_345_i17_3_lut_4_lut (.A(n11778), .B(n22242), .C(in_port[3]), 
         .D(n16_adj_1333), .Z(n17_adj_569)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_345_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_349_i17_3_lut_4_lut (.A(n11778), .B(n22242), .C(in_port[4]), 
         .D(n16_adj_1334), .Z(n17_adj_567)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_349_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_353_i17_3_lut_4_lut (.A(n11778), .B(n22242), .C(in_port[5]), 
         .D(n16_adj_1335), .Z(n17_adj_565)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_353_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_357_i17_3_lut_4_lut (.A(n11778), .B(n22242), .C(in_port[6]), 
         .D(n16_adj_1336), .Z(n17_adj_562)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_357_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_574_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n11714), 
         .D(n16392), .Z(n22141)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_574_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_598_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n7762), 
         .D(n16392), .Z(n22165)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_598_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_622_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n16312), 
         .D(n16392), .Z(n22189)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_622_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_549_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n7908), 
         .D(n7876), .Z(n22116)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_549_3_lut_4_lut.init = 16'h1000;
    LUT4 PrioSelect_117_i12_3_lut_4_lut (.A(n22254), .B(n11714), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1337)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_117_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_305_i17_3_lut_4_lut (.A(n7876), .B(n22244), .C(in_port[1]), 
         .D(n16_adj_1338), .Z(n17_adj_595)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_305_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_309_i17_3_lut_4_lut (.A(n7876), .B(n22244), .C(in_port[2]), 
         .D(n16_adj_1339), .Z(n17_adj_592)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_309_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_313_i17_3_lut_4_lut (.A(n7876), .B(n22244), .C(in_port[3]), 
         .D(n16_adj_1340), .Z(n17_adj_590)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_313_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_317_i17_3_lut_4_lut (.A(n7876), .B(n22244), .C(in_port[4]), 
         .D(n16_adj_1341), .Z(n17_adj_588)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_317_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_125 (.A(instruction[12]), .B(Z_N_377), .Z(n29)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_2_lut_adj_125.init = 16'h8888;
    LUT4 i8206_3_lut (.A(st[0]), .B(rst_n_in), .C(n1124), .Z(n3[0])) /* synthesis lut_function=(A (B (C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam i8206_3_lut.init = 16'h8484;
    LUT4 PrioSelect_121_i12_3_lut_4_lut (.A(n22254), .B(n11714), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1342)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_121_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_125_i12_3_lut_4_lut (.A(n22254), .B(n11714), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1343)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_125_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_321_i17_3_lut_4_lut (.A(n7876), .B(n22244), .C(in_port[5]), 
         .D(n16_adj_1344), .Z(n17_adj_585)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_321_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_580_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n11714), 
         .D(n7876), .Z(n22147)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_580_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_604_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n7762), 
         .D(n7876), .Z(n22171)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_604_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_628_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n16312), 
         .D(n7876), .Z(n22195)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_628_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_610_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n16312), 
         .D(n11778), .Z(n22177)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_610_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_586_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n7762), 
         .D(n11778), .Z(n22153)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_586_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_646_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n7908), 
         .D(n11778), .Z(n22213)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_646_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_568_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n11714), 
         .D(n7726), .Z(n22135)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_568_3_lut_4_lut.init = 16'h0100;
    LUT4 PrioSelect_325_i17_3_lut_4_lut (.A(n7876), .B(n22244), .C(in_port[6]), 
         .D(n16_adj_1345), .Z(n17_adj_582)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_325_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_592_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n7762), 
         .D(n7726), .Z(n22159)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_592_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_616_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n16312), 
         .D(n7726), .Z(n22183)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_616_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_652_3_lut_4_lut (.A(n10_adj_586), .B(n22277), .C(n7908), 
         .D(n7726), .Z(n22219)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_652_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_4_lut_adj_126 (.A(n19961), .B(n11804), .C(n30), .D(st_zc[4]), 
         .Z(n7696)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_4_lut_adj_126.init = 16'hc088;
    LUT4 PrioSelect_129_i12_3_lut_4_lut (.A(n22254), .B(n11714), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1346)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_129_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17159_3_lut (.A(n10_adj_596), .B(n14_adj_658), .C(n16701), .Z(n15_adj_943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17159_3_lut.init = 16'hcaca;
    LUT4 i17161_3_lut (.A(n10_adj_1347), .B(n14_adj_532), .C(n16701), 
         .Z(n15_adj_933)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17161_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_277_i17_3_lut_4_lut (.A(n16392), .B(n22244), .C(in_port[2]), 
         .D(n16_adj_1348), .Z(n17_adj_611)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_277_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i17163_3_lut (.A(n10_adj_1349), .B(n14_adj_626), .C(n16701), 
         .Z(n15_adj_924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17163_3_lut.init = 16'hcaca;
    LUT4 i17165_3_lut (.A(n10_adj_1350), .B(n14_adj_656), .C(n16701), 
         .Z(n15_adj_916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17165_3_lut.init = 16'hcaca;
    LUT4 i17167_3_lut (.A(n10_adj_1351), .B(n14_adj_660), .C(n16701), 
         .Z(n15_adj_903)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17167_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_273_i17_3_lut_4_lut (.A(n16392), .B(n22244), .C(in_port[1]), 
         .D(n16_adj_1352), .Z(n17_adj_613)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_273_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_133_i12_3_lut_4_lut (.A(n22254), .B(n11714), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1353)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_133_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_281_i17_3_lut_4_lut (.A(n16392), .B(n22244), .C(in_port[3]), 
         .D(n16_adj_1354), .Z(n17_adj_608)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_281_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_285_i17_3_lut_4_lut (.A(n16392), .B(n22244), .C(in_port[4]), 
         .D(n16_adj_1355), .Z(n17_adj_606)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_285_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i17169_3_lut (.A(n10_adj_1042), .B(n14_adj_662), .C(n16701), 
         .Z(n15_adj_889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17169_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_289_i17_3_lut_4_lut (.A(n16392), .B(n22244), .C(in_port[5]), 
         .D(n16_adj_1356), .Z(n17_adj_604)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_289_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_293_i17_3_lut_4_lut (.A(n16392), .B(n22244), .C(in_port[6]), 
         .D(n16_adj_1357), .Z(n17_adj_601)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_293_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_241_i17_3_lut_4_lut (.A(n7726), .B(n22244), .C(in_port[1]), 
         .D(n16_adj_1358), .Z(n17_adj_638)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_241_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_245_i17_3_lut_4_lut (.A(n7726), .B(n22244), .C(in_port[2]), 
         .D(n16_adj_1359), .Z(n17_adj_636)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_245_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_201_i19_4_lut (.A(n17_adj_1360), .B(in_port[7]), .C(n22103), 
         .D(n346[3]), .Z(n523)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_201_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_109_i15_3_lut_4_lut (.A(n22254), .B(n11714), .C(n1108[0]), 
         .D(n5_adj_1148), .Z(n15_adj_1181)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_109_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_205_i19_4_lut (.A(n17_adj_1361), .B(in_port[0]), .C(n22206), 
         .D(n346[4]), .Z(n527)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_205_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_249_i17_3_lut_4_lut (.A(n7726), .B(n22244), .C(in_port[3]), 
         .D(n16_adj_1362), .Z(n17_adj_634)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_249_i17_3_lut_4_lut.init = 16'hf780;
    CCU2D add_21_11 (.A0(address[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(address[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14269), .COUT(n14270), .S0(n18[9]), .S1(n18[10]));   // f:/home/mini-mcu/step_fpga/mcu.v(217[27:35])
    defparam add_21_11.INIT0 = 16'h5aaa;
    defparam add_21_11.INIT1 = 16'h5aaa;
    defparam add_21_11.INJECT1_0 = "NO";
    defparam add_21_11.INJECT1_1 = "NO";
    LUT4 PrioSelect_253_i17_3_lut_4_lut (.A(n7726), .B(n22244), .C(in_port[4]), 
         .D(n16_adj_1363), .Z(n17_adj_630)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_253_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_127 (.A(instruction[10]), .B(instruction[11]), .Z(n7762)) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam i1_2_lut_adj_127.init = 16'h2222;
    LUT4 PrioSelect_257_i17_3_lut_4_lut (.A(n7726), .B(n22244), .C(in_port[5]), 
         .D(n16_adj_1364), .Z(n17_adj_628)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_257_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_261_i17_3_lut_4_lut (.A(n7726), .B(n22244), .C(in_port[6]), 
         .D(n16_adj_1365), .Z(n17_adj_622)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam PrioSelect_261_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_137_i15_3_lut_4_lut (.A(n22254), .B(n11714), .C(n1108[7]), 
         .D(n9_adj_777), .Z(n15_adj_841)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_137_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_233_i19_4_lut (.A(n17_adj_1366), .B(in_port[7]), .C(n22206), 
         .D(n346[4]), .Z(n555)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_233_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_237_i19_4_lut (.A(n17_adj_1367), .B(in_port[0]), .C(n22204), 
         .D(n346[5]), .Z(n559)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_237_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_265_i19_4_lut (.A(n17_adj_1368), .B(in_port[7]), .C(n22204), 
         .D(n346[5]), .Z(n596)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_265_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_269_i19_4_lut (.A(n17_adj_1369), .B(in_port[0]), .C(n22203), 
         .D(n346[6]), .Z(n600)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_269_i19_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_adj_128 (.A(n7762), .B(n15_adj_833), .C(n16590), .D(n22280), 
         .Z(clk_in_c_enable_52)) /* synthesis lut_function=(A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut_adj_128.init = 16'h8a88;
    LUT4 i13423_4_lut (.A(n22279), .B(n22243), .C(n22270), .D(n22273), 
         .Z(n16590)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i13423_4_lut.init = 16'h8000;
    LUT4 PrioSelect_297_i19_4_lut (.A(n17_adj_1370), .B(in_port[7]), .C(n22203), 
         .D(n346[6]), .Z(n628)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_297_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_137_i10_3_lut_4_lut (.A(n22259), .B(n11714), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1371)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_137_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_301_i19_4_lut (.A(n17_adj_1372), .B(in_port[0]), .C(n22202), 
         .D(n346[7]), .Z(n632)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_301_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_329_i19_4_lut (.A(n17_adj_1373), .B(in_port[7]), .C(n22202), 
         .D(n346[7]), .Z(n661)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_329_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_333_i19_4_lut (.A(n17_adj_1374), .B(in_port[0]), .C(n22201), 
         .D(n346[8]), .Z(n665)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_333_i19_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_rep_693_3_lut_4_lut (.A(n8050), .B(n10_adj_586), .C(n9_adj_707), 
         .D(n8_adj_708), .Z(n22260)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;
    defparam i1_2_lut_rep_693_3_lut_4_lut.init = 16'heee0;
    LUT4 i1_2_lut_adj_129 (.A(instruction[11]), .B(instruction[10]), .Z(n16312)) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i1_2_lut_adj_129.init = 16'h2222;
    LUT4 i6_3_lut_4_lut (.A(n8_adj_708), .B(n10_adj_698), .C(n22278), 
         .D(n4), .Z(n16_adj_1375)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(383[17:25])
    defparam i6_3_lut_4_lut.init = 16'he000;
    LUT4 i13383_2_lut_rep_676_3_lut (.A(n8_adj_708), .B(n10_adj_698), .C(n11916), 
         .Z(n22243)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(383[17:25])
    defparam i13383_2_lut_rep_676_3_lut.init = 16'he0e0;
    LUT4 i13409_3_lut_4_lut_4_lut (.A(n8_adj_708), .B(n10_adj_698), .C(n22325), 
         .D(n9_adj_707), .Z(n16574)) /* synthesis lut_function=(A (C)+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(383[17:25])
    defparam i13409_3_lut_4_lut_4_lut.init = 16'he0a0;
    LUT4 PrioSelect_361_i19_4_lut (.A(n17_adj_1376), .B(in_port[7]), .C(n22201), 
         .D(n346[8]), .Z(n693)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_361_i19_4_lut.init = 16'hc0ca;
    LUT4 i1578_3_lut_4_lut (.A(n22259), .B(n11714), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1377)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i1578_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_365_i19_4_lut (.A(n17_adj_1378), .B(in_port[0]), .C(n22200), 
         .D(n346[9]), .Z(n697)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_365_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_393_i19_4_lut (.A(n17_adj_1379), .B(in_port[7]), .C(n22200), 
         .D(n346[9]), .Z(n734)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_393_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_133_i13_3_lut_4_lut (.A(n22259), .B(n11714), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1380)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_133_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_397_i19_4_lut (.A(n17_adj_1381), .B(in_port[0]), .C(n22199), 
         .D(n346[10]), .Z(n738)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_397_i19_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_adj_130 (.A(n16392), .B(n16312), .C(n22261), .D(n22198), 
         .Z(clk_in_c_enable_76)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_130.init = 16'hcc80;
    LUT4 PrioSelect_425_i19_4_lut (.A(n17_adj_1382), .B(in_port[7]), .C(n22199), 
         .D(n346[10]), .Z(n766)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_425_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_209_i17_3_lut_4_lut (.A(n11778), .B(n22244), .C(in_port[1]), 
         .D(n16_adj_1383), .Z(n17_adj_668)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_209_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_129_i13_3_lut_4_lut (.A(n22259), .B(n11714), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1384)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_129_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_429_i19_4_lut (.A(n17_adj_1385), .B(in_port[0]), .C(n22197), 
         .D(n346[11]), .Z(n770)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_429_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_457_i19_4_lut (.A(n17_adj_1386), .B(in_port[7]), .C(n22197), 
         .D(n346[11]), .Z(n798)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_457_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_125_i13_3_lut_4_lut (.A(n22259), .B(n11714), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1387)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_125_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_461_i19_4_lut (.A(n17_adj_1388), .B(in_port[0]), .C(n22209), 
         .D(n346[12]), .Z(n802)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_461_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_489_i19_4_lut (.A(n17_adj_1389), .B(in_port[7]), .C(n22209), 
         .D(n346[12]), .Z(n830)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_489_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_121_i13_3_lut_4_lut (.A(n22259), .B(n11714), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1390)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_121_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_493_i19_4_lut (.A(n17_adj_1391), .B(in_port[0]), .C(n22256), 
         .D(n346[13]), .Z(n834)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_493_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_137_i8_4_lut (.A(n6_adj_694), .B(n7_adj_473), .C(n16282), 
         .D(n16289), .Z(n8_adj_845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_137_i8_4_lut.init = 16'hcfca;
    LUT4 PrioSelect_213_i17_3_lut_4_lut (.A(n11778), .B(n22244), .C(in_port[2]), 
         .D(n16_adj_1392), .Z(n17_adj_666)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_213_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_521_i19_4_lut (.A(n17_adj_1393), .B(in_port[7]), .C(n22256), 
         .D(n346[13]), .Z(n862)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_521_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_117_i13_3_lut_4_lut (.A(n22259), .B(n11714), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1394)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_117_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_525_i19_4_lut (.A(n17_adj_1395), .B(in_port[0]), .C(n22196), 
         .D(n346[14]), .Z(n866)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_525_i19_4_lut.init = 16'hc0ca;
    LUT4 i8566_4_lut (.A(n21644), .B(rst_n_in), .C(st[2]), .D(n1124), 
         .Z(n3[2])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam i8566_4_lut.init = 16'hc088;
    LUT4 PrioSelect_113_i13_3_lut_4_lut (.A(n22259), .B(n11714), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1396)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_113_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_553_i19_4_lut (.A(n17_adj_1397), .B(in_port[7]), .C(n22196), 
         .D(n346[14]), .Z(n894)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_553_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_557_i19_4_lut (.A(n17_adj_1398), .B(in_port[0]), .C(n22241), 
         .D(n346[15]), .Z(n898)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_557_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_585_i19_4_lut (.A(n17_adj_1399), .B(in_port[7]), .C(n22241), 
         .D(n346[15]), .Z(n926)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_585_i19_4_lut.init = 16'hc0ca;
    LUT4 mux_628_i6_3_lut (.A(n18[5]), .B(address[5]), .C(clk_in_c_enable_109), 
         .Z(n1844[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i6_3_lut.init = 16'hacac;
    LUT4 i1_4_lut_adj_131 (.A(instruction[12]), .B(n16364), .C(instruction[14]), 
         .D(instruction[17]), .Z(out_port_7__N_232)) /* synthesis lut_function=(A (B (C (D)))+!A (B (C (D)+!C !(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i1_4_lut_adj_131.init = 16'hc004;
    LUT4 PrioSelect_113_i14_3_lut_4_lut (.A(n22257), .B(n11714), .C(Z_N_387[1]), 
         .D(n13_adj_1396), .Z(n14_adj_757)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_113_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_117_i14_3_lut_4_lut (.A(n22257), .B(n11714), .C(Z_N_387[2]), 
         .D(n13_adj_1394), .Z(n14_adj_773)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_117_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_217_i17_3_lut_4_lut (.A(n11778), .B(n22244), .C(in_port[3]), 
         .D(n16_adj_1400), .Z(n17_adj_651)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_217_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i6954_1_lut (.A(out_port_7__N_232), .Z(n10012)) /* synthesis lut_function=(!(A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i6954_1_lut.init = 16'h5555;
    LUT4 PrioSelect_121_i14_3_lut_4_lut (.A(n22257), .B(n11714), .C(Z_N_387[3]), 
         .D(n13_adj_1390), .Z(n14_adj_767)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_121_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_221_i17_3_lut_4_lut (.A(n11778), .B(n22244), .C(in_port[4]), 
         .D(n16_adj_1401), .Z(n17_adj_647)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_221_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_125_i14_3_lut_4_lut (.A(n22257), .B(n11714), .C(Z_N_387[4]), 
         .D(n13_adj_1387), .Z(n14_adj_760)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_125_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut (.A(instruction[13]), .B(instruction[16]), .C(instruction[15]), 
         .Z(n16364)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i1_3_lut.init = 16'h1010;
    LUT4 Mux_6_i15_3_lut (.A(n7_adj_462), .B(n14_adj_463), .C(instruction[11]), 
         .Z(s_N_294[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_6_i15_3_lut.init = 16'hcaca;
    LUT4 Mux_5_i15_3_lut (.A(n7_adj_609), .B(n14_adj_705), .C(instruction[11]), 
         .Z(s_N_294[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 Mux_5_i14_3_lut (.A(n19766), .B(n13_adj_744), .C(instruction[10]), 
         .Z(n14_adj_705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_5_i14_3_lut.init = 16'hcaca;
    LUT4 Mux_4_i15_3_lut (.A(n7_adj_476), .B(n14_adj_709), .C(instruction[11]), 
         .Z(s_N_294[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_4_i15_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_225_i17_3_lut_4_lut (.A(n11778), .B(n22244), .C(in_port[5]), 
         .D(n16_adj_1402), .Z(n17_adj_645)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_225_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_129_i14_3_lut_4_lut (.A(n22257), .B(n11714), .C(Z_N_387[5]), 
         .D(n13_adj_1384), .Z(n14_adj_770)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_129_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 Mux_4_i14_3_lut (.A(n19760), .B(n13_adj_515), .C(instruction[10]), 
         .Z(n14_adj_709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[48:57])
    defparam Mux_4_i14_3_lut.init = 16'hcaca;
    LUT4 i17586_4_lut (.A(n22120), .B(n22122), .C(n22121), .D(n213[14]), 
         .Z(n19390)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17586_4_lut.init = 16'haaab;
    LUT4 i1_3_lut_adj_132 (.A(instruction[14]), .B(n16364), .C(instruction[17]), 
         .Z(port_id_7__N_215)) /* synthesis lut_function=(A (B (C))+!A !((C)+!B)) */ ;
    defparam i1_3_lut_adj_132.init = 16'h8484;
    LUT4 i6952_1_lut (.A(port_id_7__N_215), .Z(n10010)) /* synthesis lut_function=(!(A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i6952_1_lut.init = 16'h5555;
    LUT4 i47_3_lut (.A(port_id_7__N_200[1]), .B(instruction[1]), .C(instruction[12]), 
         .Z(n23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i47_3_lut.init = 16'hcaca;
    LUT4 i16495_3_lut (.A(n19663), .B(n19664), .C(instruction[7]), .Z(port_id_7__N_200[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16495_3_lut.init = 16'hcaca;
    LUT4 i47_3_lut_adj_133 (.A(port_id_7__N_200[2]), .B(instruction[2]), 
         .C(instruction[12]), .Z(n23_adj_485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i47_3_lut_adj_133.init = 16'hcaca;
    LUT4 i16450_3_lut (.A(n19618), .B(n19619), .C(instruction[7]), .Z(port_id_7__N_200[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16450_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_229_i17_3_lut_4_lut (.A(n11778), .B(n22244), .C(in_port[6]), 
         .D(n16_adj_1403), .Z(n17_adj_643)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_229_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i47_3_lut_adj_134 (.A(port_id_7__N_200[3]), .B(instruction[3]), 
         .C(instruction[12]), .Z(n23_adj_486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i47_3_lut_adj_134.init = 16'hcaca;
    LUT4 i16420_3_lut (.A(n19588), .B(n19589), .C(instruction[7]), .Z(port_id_7__N_200[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16420_3_lut.init = 16'hcaca;
    LUT4 i47_3_lut_adj_135 (.A(port_id_7__N_200[4]), .B(instruction[4]), 
         .C(instruction[12]), .Z(n23_adj_487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i47_3_lut_adj_135.init = 16'hcaca;
    LUT4 i16435_3_lut (.A(n19603), .B(n19604), .C(instruction[7]), .Z(port_id_7__N_200[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16435_3_lut.init = 16'hcaca;
    LUT4 i47_3_lut_adj_136 (.A(port_id_7__N_200[5]), .B(instruction[5]), 
         .C(instruction[12]), .Z(n23_adj_488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i47_3_lut_adj_136.init = 16'hcaca;
    LUT4 i16480_3_lut (.A(n19648), .B(n19649), .C(instruction[7]), .Z(port_id_7__N_200[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16480_3_lut.init = 16'hcaca;
    LUT4 i47_3_lut_adj_137 (.A(port_id_7__N_200[6]), .B(instruction[6]), 
         .C(instruction[12]), .Z(n23_adj_489)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i47_3_lut_adj_137.init = 16'hcaca;
    LUT4 i16614_3_lut (.A(n19782), .B(n19783), .C(instruction[7]), .Z(port_id_7__N_200[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16614_3_lut.init = 16'hcaca;
    LUT4 i47_3_lut_adj_138 (.A(port_id_7__N_200[7]), .B(instruction[7]), 
         .C(instruction[12]), .Z(n23_adj_490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i47_3_lut_adj_138.init = 16'hcaca;
    LUT4 mux_628_i5_3_lut (.A(n18[4]), .B(address[4]), .C(clk_in_c_enable_109), 
         .Z(n1844[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i5_3_lut.init = 16'hacac;
    LUT4 PrioSelect_133_i14_3_lut_4_lut (.A(n22257), .B(n11714), .C(Z_N_387[6]), 
         .D(n13_adj_1380), .Z(n14_adj_750)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_133_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_469_i11_3_lut_4_lut (.A(n22245), .B(n7908), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1404)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_469_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_109_i14_3_lut_4_lut (.A(n22257), .B(n11714), .C(Z_N_387[0]), 
         .D(n10_adj_1377), .Z(n14_adj_1180)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_109_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_465_i11_3_lut_4_lut (.A(n22245), .B(n7908), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1405)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_465_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_473_i11_3_lut_4_lut (.A(n22245), .B(n7908), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1406)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_473_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_137_i14_3_lut_4_lut (.A(n22257), .B(n11714), .C(Z_N_387[7]), 
         .D(n10_adj_1371), .Z(n14_adj_840)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_137_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17721_4_lut (.A(n22193), .B(n22195), .C(n22194), .D(n213[11]), 
         .Z(n18838)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17721_4_lut.init = 16'haaab;
    LUT4 PrioSelect_477_i11_3_lut_4_lut (.A(n22245), .B(n7908), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1407)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_477_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_628_i4_3_lut (.A(n18[3]), .B(address[3]), .C(clk_in_c_enable_109), 
         .Z(n1844[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i4_3_lut.init = 16'hacac;
    LUT4 i8511_4_lut (.A(s_11_7), .B(n16318), .C(n14_adj_709), .D(n16358), 
         .Z(n6_adj_1408)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8511_4_lut.init = 16'h3022;
    LUT4 PrioSelect_481_i11_3_lut_4_lut (.A(n22245), .B(n7908), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1409)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_481_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_485_i11_3_lut_4_lut (.A(n22245), .B(n7908), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1410)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_485_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_489_i11_3_lut_4_lut (.A(n22246), .B(n7908), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1411)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_489_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_149_i11_3_lut_4_lut (.A(n22229), .B(n11714), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1412)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_149_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_145_i11_3_lut_4_lut (.A(n22229), .B(n11714), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1413)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_145_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_153_i11_3_lut_4_lut (.A(n22229), .B(n11714), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1414)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_153_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_461_i11_3_lut_4_lut (.A(n22246), .B(n7908), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1415)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_461_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 C_N_336_0__bdd_4_lut_18216 (.A(C_N_336[0]), .B(out_port_7__N_217[0]), 
         .C(instruction[0]), .D(instruction[2]), .Z(n21790)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+(C (D))))) */ ;
    defparam C_N_336_0__bdd_4_lut_18216.init = 16'h0311;
    LUT4 i17747_4_lut (.A(n22193), .B(n22195), .C(n22194), .D(n18796), 
         .Z(n20349)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17747_4_lut.init = 16'habaa;
    LUT4 i15606_4_lut (.A(n22192), .B(n22191), .C(n22190), .D(n213[11]), 
         .Z(n18796)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15606_4_lut.init = 16'h5554;
    LUT4 mux_628_i2_3_lut (.A(n18[1]), .B(address[1]), .C(clk_in_c_enable_109), 
         .Z(n1844[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i2_3_lut.init = 16'hacac;
    LUT4 mux_628_i1_3_lut (.A(n18[0]), .B(address[0]), .C(clk_in_c_enable_109), 
         .Z(n1844[0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i1_3_lut.init = 16'hacac;
    PFUMX C_N_340_7__I_0_587_i16 (.BLUT(n8_adj_1416), .ALUT(n14_adj_1417), 
          .C0(n16636), .Z(n16_adj_843)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 mux_628_i3_3_lut (.A(n18[2]), .B(address[2]), .C(clk_in_c_enable_109), 
         .Z(n1844[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i3_3_lut.init = 16'hacac;
    LUT4 PrioSelect_157_i11_3_lut_4_lut (.A(n22229), .B(n11714), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1418)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_157_i11_3_lut_4_lut.init = 16'hfd20;
    PFUMX i106 (.BLUT(n14422), .ALUT(n77), .C0(instruction[15]), .Z(n50));
    LUT4 PrioSelect_465_i17_3_lut_4_lut (.A(n11778), .B(n22247), .C(in_port[1]), 
         .D(n16_adj_1419), .Z(n17_adj_484)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_465_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_161_i11_3_lut_4_lut (.A(n22229), .B(n11714), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1420)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_161_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17758_4_lut (.A(n22187), .B(n22189), .C(n22188), .D(n213[10]), 
         .Z(n18654)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17758_4_lut.init = 16'haaab;
    LUT4 i17491_4_lut_4_lut (.A(n22129), .B(n16800), .C(n22128), .D(n22127), 
         .Z(n16810)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i17491_4_lut_4_lut.init = 16'hffef;
    LUT4 PrioSelect_469_i17_3_lut_4_lut (.A(n11778), .B(n22247), .C(in_port[2]), 
         .D(n16_adj_1421), .Z(n17_adj_478)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_469_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_473_i17_3_lut_4_lut (.A(n11778), .B(n22247), .C(in_port[3]), 
         .D(n16_adj_1422), .Z(n17_adj_475)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_473_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i8568_4_lut (.A(n2641[3]), .B(rst_n_in), .C(st[4]), .D(n1124), 
         .Z(n3[4])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam i8568_4_lut.init = 16'hc088;
    LUT4 mux_1308_i4_4_lut (.A(stack_N_397[4]), .B(st[4]), .C(n14459), 
         .D(n8_adj_1289), .Z(n2641[3])) /* synthesis lut_function=(A (B (C+(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_1308_i4_4_lut.init = 16'haca3;
    LUT4 PrioSelect_477_i17_3_lut_4_lut (.A(n11778), .B(n22247), .C(in_port[4]), 
         .D(n16_adj_1423), .Z(n17_adj_472)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_477_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_165_i11_3_lut_4_lut (.A(n22229), .B(n11714), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1424)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_165_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_628_i12_3_lut (.A(n18[11]), .B(address[11]), .C(clk_in_c_enable_109), 
         .Z(n1844[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i12_3_lut.init = 16'hacac;
    LUT4 mux_628_i11_3_lut (.A(n18[10]), .B(address[10]), .C(clk_in_c_enable_109), 
         .Z(n1844[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i11_3_lut.init = 16'hacac;
    LUT4 i1738_3_lut_4_lut (.A(n8647), .B(n11714), .C(n7_adj_462), .D(n7_adj_481), 
         .Z(n10_adj_791)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1738_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_481_i17_3_lut_4_lut (.A(n11778), .B(n22247), .C(in_port[5]), 
         .D(n16_adj_1425), .Z(n17_adj_470)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_481_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_485_i17_3_lut_4_lut (.A(n11778), .B(n22247), .C(in_port[6]), 
         .D(n16_adj_1426), .Z(n17_adj_467)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam PrioSelect_485_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1754_3_lut_4_lut (.A(n8647), .B(n11714), .C(n7_adj_609), .D(n7_c), 
         .Z(n10_adj_787)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1754_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1770_3_lut_4_lut (.A(n8647), .B(n11714), .C(n7_adj_476), .D(n7_adj_462), 
         .Z(n10_adj_794)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1770_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1116_1_lut (.A(st[0]), .Z(stack_N_397[0])) /* synthesis lut_function=(!(A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(284[52:61])
    defparam i1116_1_lut.init = 16'h5555;
    LUT4 i17693_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22248), .B(n7908), .C(n22245), 
         .D(n22246), .Z(n19010)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17693_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h4ccc;
    LUT4 i1_2_lut_3_lut_4_lut_adj_139 (.A(n22261), .B(n22205), .C(n7876), 
         .D(n16312), .Z(clk_in_c_enable_82)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_139.init = 16'hb000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_140 (.A(n22261), .B(n22205), .C(n7726), 
         .D(n16312), .Z(clk_in_c_enable_70)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_140.init = 16'hb000;
    LUT4 PrioSelect_489_i12_3_lut_4_lut (.A(n22248), .B(n7908), .C(Z_N_378[7]), 
         .D(n11_adj_1411), .Z(n12_adj_1427)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_489_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_461_i12_3_lut_4_lut (.A(n22248), .B(n7908), .C(Z_N_378[0]), 
         .D(n11_adj_1415), .Z(n12_adj_1428)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_461_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17764_4_lut (.A(n22187), .B(n22189), .C(n22188), .D(n18612), 
         .Z(n20366)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17764_4_lut.init = 16'habaa;
    LUT4 i15422_4_lut (.A(n22186), .B(n22185), .C(n22184), .D(n213[10]), 
         .Z(n18612)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15422_4_lut.init = 16'h5554;
    LUT4 i1786_3_lut_4_lut (.A(n8647), .B(n11714), .C(n7_adj_473), .D(n7_adj_609), 
         .Z(n10_adj_779)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1786_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_205_i5_3_lut_4_lut (.A(n7762), .B(n8627), .C(n7_adj_479), 
         .D(n7_adj_473), .Z(n5_adj_1429)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_205_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i8565_4_lut (.A(n4_adj_1430), .B(rst_n_in), .C(st[1]), .D(n1124), 
         .Z(n3[1])) /* synthesis lut_function=(A (B (C))+!A (B (C (D)+!C !(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam i8565_4_lut.init = 16'hc084;
    LUT4 PrioSelect_169_i11_3_lut_4_lut (.A(n22230), .B(n11714), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1431)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_169_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_141_i11_3_lut_4_lut (.A(n22230), .B(n11714), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1432)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_141_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_521_i9_3_lut_4_lut (.A(n22093), .B(n7908), .C(n14_adj_501), 
         .D(C), .Z(n9_adj_631)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_521_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_465_i12_3_lut_4_lut (.A(n22250), .B(n7908), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1433)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_465_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_469_i12_3_lut_4_lut (.A(n22250), .B(n7908), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1434)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_469_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_473_i12_3_lut_4_lut (.A(n22250), .B(n7908), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1435)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_473_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1930_3_lut_4_lut (.A(n7762), .B(n8627), .C(n7_adj_481), .D(n7_adj_500), 
         .Z(n10_adj_824)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1930_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_581_i16 (.BLUT(n11_adj_1436), .ALUT(n12_adj_1437), 
          .C0(n19547), .Z(n16_adj_1119)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_477_i12_3_lut_4_lut (.A(n22250), .B(n7908), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1438)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_477_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1946_3_lut_4_lut (.A(n7762), .B(n8627), .C(n7_c), .D(n7_adj_479), 
         .Z(n10_adj_858)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1946_3_lut_4_lut.init = 16'hf780;
    LUT4 i17585_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22231), .B(n11714), .C(n22229), 
         .D(n22230), .Z(n17170)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17585_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3332;
    LUT4 i1962_3_lut_4_lut (.A(n7762), .B(n8627), .C(n7_adj_462), .D(n7_adj_481), 
         .Z(n10_adj_832)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1962_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_553_i9_3_lut_4_lut (.A(n22095), .B(n7908), .C(n14_adj_501), 
         .D(C), .Z(n9_adj_1175)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_553_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_141 (.A(n14459), .B(st[0]), .Z(n4_adj_1430)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_2_lut_adj_141.init = 16'h6666;
    PFUMX PrioSelect_577_i16 (.BLUT(n11_adj_1439), .ALUT(n12_adj_1440), 
          .C0(n19547), .Z(n16_adj_1117)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_adj_142 (.A(st[0]), .B(st[1]), .Z(stack_N_397[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_2_lut_adj_142.init = 16'h6666;
    LUT4 PrioSelect_481_i12_3_lut_4_lut (.A(n22250), .B(n7908), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1441)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_481_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_485_i12_3_lut_4_lut (.A(n22250), .B(n7908), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1442)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_485_i12_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_549_i16 (.BLUT(n11_adj_1443), .ALUT(n12_adj_1171), 
          .C0(n19363), .Z(n16_adj_1309)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 mux_628_i10_3_lut (.A(n18[9]), .B(address[9]), .C(clk_in_c_enable_109), 
         .Z(n1844[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i10_3_lut.init = 16'hacac;
    LUT4 mux_628_i9_3_lut (.A(n18[8]), .B(address[8]), .C(clk_in_c_enable_109), 
         .Z(n1844[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i9_3_lut.init = 16'hacac;
    LUT4 PrioSelect_169_i12_3_lut_4_lut (.A(n22231), .B(n11714), .C(Z_N_378[7]), 
         .D(n11_adj_1431), .Z(n12_adj_1444)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_169_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17492_4_lut (.A(n22181), .B(n22183), .C(n22182), .D(n213[9]), 
         .Z(n18321)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17492_4_lut.init = 16'haaab;
    PFUMX PrioSelect_545_i16 (.BLUT(n11_adj_1445), .ALUT(n12_adj_1169), 
          .C0(n19363), .Z(n16_adj_1307)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1978_3_lut_4_lut (.A(n7762), .B(n8627), .C(n7_adj_609), .D(n7_c), 
         .Z(n10_adj_827)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1978_3_lut_4_lut.init = 16'hf780;
    LUT4 i8493_4_lut (.A(s_9_7), .B(n16319), .C(n14_adj_709), .D(n16357), 
         .Z(n6_adj_1446)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8493_4_lut.init = 16'h3022;
    LUT4 PrioSelect_461_i15_3_lut_4_lut (.A(n22250), .B(n7908), .C(n1108[0]), 
         .D(n5_adj_732), .Z(n15_adj_952)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_461_i15_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_517_i16 (.BLUT(n11_adj_687), .ALUT(n12_adj_620), .C0(n19179), 
          .Z(n16_adj_1241)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_141_i12_3_lut_4_lut (.A(n22231), .B(n11714), .C(Z_N_378[0]), 
         .D(n11_adj_1432), .Z(n12_adj_1447)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_141_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_489_i15_3_lut_4_lut (.A(n22250), .B(n7908), .C(n1108[7]), 
         .D(n9_adj_1116), .Z(n15_adj_465)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_489_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17487_4_lut (.A(n22181), .B(n22183), .C(n22182), .D(n18368), 
         .Z(n20089)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17487_4_lut.init = 16'habaa;
    PFUMX PrioSelect_513_i16 (.BLUT(n11_adj_686), .ALUT(n12_adj_583), .C0(n19179), 
          .Z(n16_adj_1237)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i15178_4_lut (.A(n22180), .B(n22179), .C(n22178), .D(n213[9]), 
         .Z(n18368)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15178_4_lut.init = 16'h5554;
    LUT4 i1396_3_lut (.A(st_zc[0]), .B(st_zc[1]), .C(clk_in_c_enable_109), 
         .Z(n2755)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1396_3_lut.init = 16'h9696;
    LUT4 PrioSelect_489_i10_3_lut_4_lut (.A(n22252), .B(n7908), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1448)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_489_i10_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_485_i16 (.BLUT(n11_adj_1410), .ALUT(n12_adj_1442), 
          .C0(n18995), .Z(n16_adj_1426)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_169_i15_3_lut_4_lut (.A(n22232), .B(n11714), .C(n1108[7]), 
         .D(n9_adj_800), .Z(n15_adj_755)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_169_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 C_N_336_0__bdd_3_lut_18217 (.A(C_N_336[0]), .B(instruction[0]), 
         .C(instruction[2]), .Z(n21789)) /* synthesis lut_function=(!(A+(B (C)))) */ ;
    defparam C_N_336_0__bdd_3_lut_18217.init = 16'h1515;
    LUT4 i17525_4_lut (.A(n22175), .B(n22177), .C(n22176), .D(n213[8]), 
         .Z(n18286)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17525_4_lut.init = 16'haaab;
    LUT4 PrioSelect_141_i15_3_lut_4_lut (.A(n22232), .B(n11714), .C(n1108[0]), 
         .D(n5_adj_1198), .Z(n15_adj_979)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_141_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_165_i12_3_lut_4_lut (.A(n22232), .B(n11714), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1449)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_165_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2810_3_lut_4_lut (.A(n22252), .B(n7908), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1450)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i2810_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17542_4_lut (.A(n22175), .B(n22177), .C(n22176), .D(n18244), 
         .Z(n20144)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17542_4_lut.init = 16'habaa;
    PFUMX PrioSelect_481_i16 (.BLUT(n11_adj_1409), .ALUT(n12_adj_1441), 
          .C0(n18995), .Z(n16_adj_1425)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i15054_4_lut (.A(n22174), .B(n22173), .C(n22172), .D(n213[8]), 
         .Z(n18244)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15054_4_lut.init = 16'h5554;
    LUT4 PrioSelect_485_i13_3_lut_4_lut (.A(n22252), .B(n7908), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1451)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_485_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_481_i13_3_lut_4_lut (.A(n22252), .B(n7908), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1452)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_481_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1307_i4_4_lut (.A(st_zc[4]), .B(n22287), .C(clk_in_c_enable_109), 
         .D(n8_adj_1453), .Z(n2634[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !(B (C (D))+!B ((D)+!C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam mux_1307_i4_4_lut.init = 16'hac5c;
    LUT4 i3_3_lut (.A(rst_n_in), .B(n5_adj_964), .C(clk_in_c_enable_109), 
         .Z(n10021)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam i3_3_lut.init = 16'h0202;
    LUT4 C_N_336_0__bdd_4_lut_18225 (.A(C_N_336[0]), .B(out_port_7__N_217[0]), 
         .C(instruction[2]), .D(C), .Z(n21792)) /* synthesis lut_function=(!(A+(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam C_N_336_0__bdd_4_lut_18225.init = 16'h1015;
    PFUMX PrioSelect_453_i16 (.BLUT(n11_adj_1260), .ALUT(n12_adj_1284), 
          .C0(n18811), .Z(n16_adj_1316)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_4_lut_adj_143 (.A(jp), .B(n17_adj_1454), .C(n15_adj_1455), 
         .D(n16_adj_1375), .Z(n5_adj_964)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(192[9] 397[7])
    defparam i1_4_lut_adj_143.init = 16'heaaa;
    LUT4 i7_4_lut_adj_144 (.A(n22274), .B(n6978), .C(n22272), .D(n22275), 
         .Z(n17_adj_1454)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_144.init = 16'h8000;
    LUT4 i5_4_lut_adj_145 (.A(n11_adj_1456), .B(n22269), .C(n9_adj_1457), 
         .D(n22322), .Z(n15_adj_1455)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_145.init = 16'h8000;
    PFUMX PrioSelect_449_i16 (.BLUT(n11_adj_1264), .ALUT(n12_adj_1279), 
          .C0(n18811), .Z(n16_adj_1315)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i4_4_lut_adj_146 (.A(n7_adj_1458), .B(n21532), .C(instruction[12]), 
         .D(n21529), .Z(n11_adj_1456)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C))) */ ;
    defparam i4_4_lut_adj_146.init = 16'hcc8c;
    LUT4 i2_4_lut_adj_147 (.A(n11_adj_872), .B(instruction[12]), .C(n16487), 
         .D(n7_adj_1458), .Z(n9_adj_1457)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i2_4_lut_adj_147.init = 16'haaa8;
    LUT4 PrioSelect_477_i13_3_lut_4_lut (.A(n22252), .B(n7908), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1459)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_477_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1994_3_lut_4_lut (.A(n7762), .B(n8627), .C(n7_adj_476), .D(n7_adj_462), 
         .Z(n10_adj_836)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1994_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_473_i13_3_lut_4_lut (.A(n22252), .B(n7908), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1460)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_473_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_161_i12_3_lut_4_lut (.A(n22232), .B(n11714), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1461)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_161_i12_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_421_i16 (.BLUT(n11_adj_1225), .ALUT(n12_adj_1247), 
          .C0(n18627), .Z(n16_adj_1323)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 instruction_17__I_0_554_i7_2_lut (.A(instruction[13]), .B(instruction[14]), 
         .Z(n7_adj_1458)) /* synthesis lut_function=(A+!(B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(216[16:21])
    defparam instruction_17__I_0_554_i7_2_lut.init = 16'hbbbb;
    CCU2D sub_131_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Z_N_378[0]), .B1(C), .C1(GND_net), .D1(GND_net), .COUT(n14278), 
          .S1(n703[0]));   // f:/home/mini-mcu/step_fpga/mcu.v(281[61:73])
    defparam sub_131_add_2_1.INIT0 = 16'h0000;
    defparam sub_131_add_2_1.INIT1 = 16'h5999;
    defparam sub_131_add_2_1.INJECT1_0 = "NO";
    defparam sub_131_add_2_1.INJECT1_1 = "NO";
    LUT4 PrioSelect_469_i13_3_lut_4_lut (.A(n22252), .B(n7908), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1462)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_469_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_149_i12_3_lut_4_lut (.A(n22232), .B(n11714), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1463)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_149_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 C_N_336_0__bdd_3_lut_18224 (.A(out_port_7__N_217[0]), .B(instruction[2]), 
         .C(C), .Z(n21793)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;
    defparam C_N_336_0__bdd_3_lut_18224.init = 16'h4545;
    LUT4 i17564_4_lut (.A(n22169), .B(n22171), .C(n22170), .D(n213[7]), 
         .Z(n18102)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17564_4_lut.init = 16'haaab;
    PFUMX PrioSelect_417_i16 (.BLUT(n11_adj_1224), .ALUT(n12_adj_1246), 
          .C0(n18627), .Z(n16_adj_1322)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i8475_4_lut (.A(s_7_7), .B(n114), .C(n7_adj_476), .D(n7094), 
         .Z(n6_adj_1464)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8475_4_lut.init = 16'h3022;
    LUT4 PrioSelect_157_i12_3_lut_4_lut (.A(n22232), .B(n11714), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1465)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_157_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17660_4_lut (.A(n22214), .B(n22219), .C(n22218), .D(n213[13]), 
         .Z(n19206)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17660_4_lut.init = 16'haaab;
    PFUMX PrioSelect_389_i16 (.BLUT(n11_adj_1192), .ALUT(n12_adj_1205), 
          .C0(n18363), .Z(n16_adj_1329)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i2010_3_lut_4_lut (.A(n7762), .B(n8627), .C(n7_adj_473), .D(n7_adj_609), 
         .Z(n10_adj_822)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2010_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_585_i9_3_lut_4_lut (.A(n22097), .B(n7908), .C(n14_adj_501), 
         .D(C), .Z(n9_adj_1466)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam PrioSelect_585_i9_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_385_i16 (.BLUT(n11_adj_1191), .ALUT(n12_adj_1204), 
          .C0(n18363), .Z(n16_adj_1328)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_145_i12_3_lut_4_lut (.A(n22232), .B(n11714), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1467)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_145_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_153_i12_3_lut_4_lut (.A(n22232), .B(n11714), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1468)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_153_i12_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_357_i16 (.BLUT(n11_adj_1141), .ALUT(n12_adj_1154), 
          .C0(n18259), .Z(n16_adj_1336)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i3_4_lut (.A(instruction[12]), .B(n22319), .C(instruction[17]), 
         .D(n16409), .Z(n1339)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_adj_148 (.A(instruction[16]), .B(n16409), .C(n105), 
         .D(n22328), .Z(n1341)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_148.init = 16'hc4c0;
    LUT4 PrioSelect_465_i13_3_lut_4_lut (.A(n22252), .B(n7908), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1469)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_465_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_169_i10_3_lut_4_lut (.A(n22233), .B(n11714), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1470)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_169_i10_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_353_i16 (.BLUT(n11_adj_1140), .ALUT(n12_adj_1153), 
          .C0(n18259), .Z(n16_adj_1335)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17575_4_lut (.A(n22169), .B(n22171), .C(n22170), .D(n18060), 
         .Z(n20177)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17575_4_lut.init = 16'habaa;
    LUT4 i1_4_lut_4_lut_adj_149 (.A(n16392), .B(clk_in_c_enable_174), .C(n22106), 
         .D(n22222), .Z(clk_in_c_enable_28)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))) */ ;
    defparam i1_4_lut_4_lut_adj_149.init = 16'haa08;
    LUT4 i14870_4_lut (.A(n22168), .B(n22167), .C(n22166), .D(n213[7]), 
         .Z(n18060)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14870_4_lut.init = 16'h5554;
    LUT4 PrioSelect_465_i14_3_lut_4_lut (.A(n22251), .B(n7908), .C(Z_N_387[1]), 
         .D(n13_adj_1469), .Z(n14_adj_1053)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_465_i14_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_325_i16 (.BLUT(n11_adj_1029), .ALUT(n12_adj_1075), 
          .C0(n18075), .Z(n16_adj_1345)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_469_i14_3_lut_4_lut (.A(n22251), .B(n7908), .C(Z_N_387[2]), 
         .D(n13_adj_1462), .Z(n14_adj_1057)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_469_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i2_4_lut_adj_150 (.A(n14413), .B(C), .C(n75), .D(n71), .Z(C_N_304)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i2_4_lut_adj_150.init = 16'hfefa;
    LUT4 i1_2_lut_2_lut_adj_151 (.A(n16122), .B(n160), .Z(n7628)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut_adj_151.init = 16'h4444;
    LUT4 i1_4_lut_adj_152 (.A(instruction[17]), .B(n14425), .C(instruction[16]), 
         .D(n53), .Z(n75)) /* synthesis lut_function=(!(A+!(B+(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_4_lut_adj_152.init = 16'h5444;
    LUT4 i2_3_lut_3_lut_adj_153 (.A(n16122), .B(n103), .C(n160), .Z(n16239)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i2_3_lut_3_lut_adj_153.init = 16'h4040;
    LUT4 PrioSelect_473_i14_3_lut_4_lut (.A(n22251), .B(n7908), .C(Z_N_387[3]), 
         .D(n13_adj_1460), .Z(n14_adj_1055)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_473_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i108_4_lut (.A(C), .B(C_N_352[0]), .C(instruction[17]), .D(n16389), 
         .Z(n56)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i108_4_lut.init = 16'hca0a;
    LUT4 Mux_5_i31_4_lut (.A(n19946), .B(n22), .C(st_zc[4]), .D(st_zc[3]), 
         .Z(C_N_352[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(376[91:109])
    defparam Mux_5_i31_4_lut.init = 16'h0aca;
    LUT4 Mux_5_i22_4_lut (.A(n19931), .B(stack_zc_d0_20_0), .C(st_zc[2]), 
         .D(n22298), .Z(n22)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(376[91:109])
    defparam Mux_5_i22_4_lut.init = 16'h0aca;
    PFUMX PrioSelect_321_i16 (.BLUT(n11_adj_1028), .ALUT(n12_adj_1074), 
          .C0(n18075), .Z(n16_adj_1344)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i2_3_lut_adj_154 (.A(instruction[13]), .B(instruction[12]), .C(n50), 
         .Z(n14425)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i2_3_lut_adj_154.init = 16'h4040;
    LUT4 i1_2_lut_adj_155 (.A(instruction[12]), .B(instruction[15]), .Z(n16389)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_2_lut_adj_155.init = 16'h8888;
    LUT4 i1690_3_lut_4_lut (.A(n22233), .B(n11714), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1471)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i1690_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_293_i16 (.BLUT(n11_adj_766), .ALUT(n12_adj_893), .C0(n17891), 
          .Z(n16_adj_1357)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_85_i11_3_lut_4_lut_4_lut (.A(n11714), .B(port_id_7__N_200[2]), 
         .C(instruction[2]), .D(n22245), .Z(n11_adj_1472)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_85_i11_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_165_i13_3_lut_4_lut (.A(n22233), .B(n11714), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1473)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_165_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_161_i13_3_lut_4_lut (.A(n22233), .B(n11714), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1474)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_161_i13_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_289_i16 (.BLUT(n11_adj_765), .ALUT(n12_adj_896), .C0(n17891), 
          .Z(n16_adj_1356)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17537_3_lut_3_lut_4_lut_4_lut (.A(n11714), .B(n22124), .C(n22125), 
         .D(n22245), .Z(n16802)) /* synthesis lut_function=(A ((C)+!B)+!A ((C+!(D))+!B)) */ ;
    defparam i17537_3_lut_3_lut_4_lut_4_lut.init = 16'hf3f7;
    LUT4 i1_4_lut_adj_156 (.A(n48), .B(n66), .C(n6_adj_1475), .D(n11196), 
         .Z(n71)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_4_lut_adj_156.init = 16'hfeff;
    LUT4 i2_4_lut_adj_157 (.A(instruction[15]), .B(instruction[12]), .C(n5_adj_861), 
         .D(instruction[14]), .Z(n6_adj_1475)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B (C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i2_4_lut_adj_157.init = 16'h7673;
    PFUMX PrioSelect_261_i16 (.BLUT(n11_adj_1476), .ALUT(n12_adj_1477), 
          .C0(n17707), .Z(n16_adj_1365)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i8146_3_lut (.A(instruction[16]), .B(instruction[15]), .C(instruction[13]), 
         .Z(n11196)) /* synthesis lut_function=(A+!(B (C)+!B !(C))) */ ;
    defparam i8146_3_lut.init = 16'hbebe;
    LUT4 PrioSelect_81_i11_3_lut_4_lut_4_lut (.A(n11714), .B(port_id_7__N_200[1]), 
         .C(instruction[1]), .D(n22245), .Z(n11_adj_1478)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_81_i11_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_97_i11_3_lut_4_lut_4_lut (.A(n11714), .B(port_id_7__N_200[5]), 
         .C(instruction[5]), .D(n22245), .Z(n11_adj_1479)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_97_i11_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX PrioSelect_257_i16 (.BLUT(n11_adj_1480), .ALUT(n12_adj_1481), 
          .C0(n17707), .Z(n16_adj_1364)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_101_i11_3_lut_4_lut_4_lut (.A(n11714), .B(port_id_7__N_200[6]), 
         .C(instruction[6]), .D(n22245), .Z(n11_adj_1482)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_101_i11_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_477_i14_3_lut_4_lut (.A(n22251), .B(n7908), .C(Z_N_387[4]), 
         .D(n13_adj_1459), .Z(n14_adj_1054)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_477_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_89_i11_3_lut_4_lut_4_lut (.A(n11714), .B(port_id_7__N_200[3]), 
         .C(instruction[3]), .D(n22245), .Z(n11_adj_1483)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_89_i11_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_481_i14_3_lut_4_lut (.A(n22251), .B(n7908), .C(Z_N_387[5]), 
         .D(n13_adj_1452), .Z(n14_adj_1056)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_481_i14_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_229_i16 (.BLUT(n11_adj_1484), .ALUT(n12_adj_1485), 
          .C0(n17523), .Z(n16_adj_1403)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_157_i13_3_lut_4_lut (.A(n22233), .B(n11714), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1486)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_157_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_153_i13_3_lut_4_lut (.A(n22233), .B(n11714), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1487)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_153_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_149_i13_3_lut_4_lut (.A(n22233), .B(n11714), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1488)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_149_i13_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_225_i16 (.BLUT(n11_adj_1489), .ALUT(n12_adj_1490), 
          .C0(n17523), .Z(n16_adj_1402)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i2_4_lut_adj_158 (.A(n14423), .B(Z), .C(n83_adj_1491), .D(n71), 
         .Z(Z_N_356)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i2_4_lut_adj_158.init = 16'hfefa;
    LUT4 i2_3_lut_adj_159 (.A(instruction[13]), .B(instruction[17]), .C(n64_adj_1492), 
         .Z(n14423)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i2_3_lut_adj_159.init = 16'h1010;
    PFUMX PrioSelect_197_i16 (.BLUT(n11_adj_673), .ALUT(n12_adj_1493), .C0(n17339), 
          .Z(n16_adj_1494)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_4_lut_adj_160 (.A(instruction[12]), .B(n16236), .C(n14417), 
         .D(n8070), .Z(n83_adj_1491)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i1_4_lut_adj_160.init = 16'ha0a8;
    LUT4 i8_4_lut_adj_161 (.A(n16532), .B(n16596), .C(n55), .D(Z_N_387[1]), 
         .Z(n16236)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i8_4_lut_adj_161.init = 16'h0010;
    PFUMX PrioSelect_193_i16 (.BLUT(n11_adj_672), .ALUT(n12_adj_1495), .C0(n17339), 
          .Z(n16_adj_1496)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_93_i11_3_lut_4_lut_4_lut (.A(n11714), .B(port_id_7__N_200[4]), 
         .C(instruction[4]), .D(n22245), .Z(n11_adj_1497)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_93_i11_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 i2_3_lut_adj_162 (.A(instruction[15]), .B(instruction[14]), .C(n61), 
         .Z(n14417)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(214[13] 386[20])
    defparam i2_3_lut_adj_162.init = 16'h2020;
    LUT4 i13428_4_lut (.A(Z_N_387[2]), .B(Z_N_387[3]), .C(Z_N_387[6]), 
         .D(n16508), .Z(n16596)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13428_4_lut.init = 16'hfffe;
    LUT4 and_168_i3_2_lut (.A(s_N_294[2]), .B(instruction[2]), .Z(Z_N_387[2])) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(351[112:121])
    defparam and_168_i3_2_lut.init = 16'h8888;
    LUT4 and_168_i4_2_lut (.A(s_N_294[3]), .B(instruction[3]), .Z(Z_N_387[3])) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(351[112:121])
    defparam and_168_i4_2_lut.init = 16'h8888;
    PFUMX PrioSelect_165_i16 (.BLUT(n11_adj_1424), .ALUT(n12_adj_1449), 
          .C0(n17155), .Z(n16_adj_1498)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 and_168_i7_2_lut (.A(s_N_294[6]), .B(instruction[6]), .Z(Z_N_387[6])) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(351[112:121])
    defparam and_168_i7_2_lut.init = 16'h8888;
    LUT4 and_168_i1_2_lut (.A(out_port_7__N_217[0]), .B(instruction[0]), 
         .Z(Z_N_387[0])) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(351[112:121])
    defparam and_168_i1_2_lut.init = 16'h8888;
    PFUMX PrioSelect_161_i16 (.BLUT(n11_adj_1420), .ALUT(n12_adj_1461), 
          .C0(n17155), .Z(n16_adj_1499)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 and_168_i2_2_lut (.A(s_N_294[1]), .B(instruction[1]), .Z(Z_N_387[1])) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(351[112:121])
    defparam and_168_i2_2_lut.init = 16'h8888;
    LUT4 and_168_i5_2_lut (.A(s_N_294[4]), .B(instruction[4]), .Z(Z_N_387[4])) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(351[112:121])
    defparam and_168_i5_2_lut.init = 16'h8888;
    LUT4 and_168_i6_2_lut (.A(s_N_294[5]), .B(instruction[5]), .Z(Z_N_387[5])) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(351[112:121])
    defparam and_168_i6_2_lut.init = 16'h8888;
    PFUMX PrioSelect_133_i16 (.BLUT(n11_adj_1296), .ALUT(n12_adj_1353), 
          .C0(n16971), .Z(n16_adj_1500)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_485_i14_3_lut_4_lut (.A(n22251), .B(n7908), .C(Z_N_387[6]), 
         .D(n13_adj_1451), .Z(n14_adj_1051)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_485_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i47_3_lut_adj_163 (.A(port_id_7__N_200[0]), .B(instruction[0]), 
         .C(instruction[12]), .Z(n23_adj_593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(404[5] 423[12])
    defparam i47_3_lut_adj_163.init = 16'hcaca;
    PFUMX PrioSelect_129_i16 (.BLUT(n11_adj_1286), .ALUT(n12_adj_1346), 
          .C0(n16971), .Z(n16_adj_1501)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i16510_3_lut (.A(n19678), .B(n19679), .C(instruction[7]), .Z(port_id_7__N_200[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16510_3_lut.init = 16'hcaca;
    LUT4 PrioSelect_145_i13_3_lut_4_lut (.A(n22233), .B(n11714), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1502)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_145_i13_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_101_i16 (.BLUT(n11_adj_1482), .ALUT(n12_adj_1503), 
          .C0(n16727), .Z(n16_adj_1275)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17344_3_lut_4_lut (.A(n22219), .B(n22102), .C(n14_adj_1504), 
         .D(n10_adj_1269), .Z(n15_adj_1505)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17344_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i18405 (.BLUT(n22308), .ALUT(n22309), .C0(instruction[16]), 
          .Z(n11916));
    LUT4 i17334_3_lut_4_lut (.A(n22219), .B(n22102), .C(n14_adj_1506), 
         .D(n10_adj_1257), .Z(n15_adj_460)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17334_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n22222), 
         .C(n7876), .D(n22106), .Z(clk_in_c_enable_34)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hc0e0;
    LUT4 i17628_4_lut (.A(n22163), .B(n22165), .C(n22164), .D(n213[6]), 
         .Z(n17918)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17628_4_lut.init = 16'haaab;
    PFUMX PrioSelect_97_i16 (.BLUT(n11_adj_1479), .ALUT(n12_adj_1507), .C0(n16727), 
          .Z(n16_adj_1274)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_145_i14_3_lut_4_lut (.A(n22234), .B(n11714), .C(Z_N_387[1]), 
         .D(n13_adj_1502), .Z(n14_adj_783)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_145_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_628_i8_3_lut (.A(n18[7]), .B(address[7]), .C(clk_in_c_enable_109), 
         .Z(n1844[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i8_3_lut.init = 16'hacac;
    LUT4 PrioSelect_461_i14_3_lut_4_lut (.A(n22251), .B(n7908), .C(Z_N_387[0]), 
         .D(n10_adj_1450), .Z(n14_adj_951)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_461_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_105_i12_3_lut_4_lut_4_lut (.A(n11714), .B(n11_adj_1218), 
         .C(Z_N_378[7]), .D(n22248), .Z(n12_adj_1508)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_105_i12_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 i17656_4_lut (.A(n22163), .B(n22165), .C(n22164), .D(n17876), 
         .Z(n20258)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17656_4_lut.init = 16'habaa;
    LUT4 i14686_4_lut (.A(n22162), .B(n22161), .C(n22160), .D(n213[6]), 
         .Z(n17876)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14686_4_lut.init = 16'h5554;
    LUT4 PrioSelect_149_i14_3_lut_4_lut (.A(n22234), .B(n11714), .C(Z_N_387[2]), 
         .D(n13_adj_1488), .Z(n14_adj_797)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_149_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17548_3_lut_3_lut_4_lut_4_lut (.A(n11714), .B(n22128), .C(n22129), 
         .D(n22248), .Z(n16701)) /* synthesis lut_function=(A ((C)+!B)+!A ((C+!(D))+!B)) */ ;
    defparam i17548_3_lut_3_lut_4_lut_4_lut.init = 16'hf3f7;
    PFUMX mux_334_i2 (.BLUT(n1742[1]), .ALUT(n1194[1]), .C0(n1341), .Z(n1238[1]));
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_164 (.A(clk_in_c_enable_174), .B(n22222), 
         .C(n7726), .D(n22106), .Z(clk_in_c_enable_22)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_164.init = 16'hc0e0;
    PFUMX mux_334_i3 (.BLUT(n1742[2]), .ALUT(n1194[2]), .C0(n1341), .Z(n1238[2]));
    LUT4 mux_628_i7_3_lut (.A(n18[6]), .B(address[6]), .C(clk_in_c_enable_109), 
         .Z(n1844[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[17:28])
    defparam mux_628_i7_3_lut.init = 16'hacac;
    LUT4 PrioSelect_489_i14_3_lut_4_lut (.A(n22251), .B(n7908), .C(Z_N_387[7]), 
         .D(n10_adj_1448), .Z(n14_adj_464)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_489_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_153_i14_3_lut_4_lut (.A(n22234), .B(n11714), .C(Z_N_387[3]), 
         .D(n13_adj_1487), .Z(n14_adj_790)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_153_i14_3_lut_4_lut.init = 16'hfd20;
    PFUMX mux_334_i4 (.BLUT(n1742[3]), .ALUT(n1194[3]), .C0(n1341), .Z(n1238[3]));
    LUT4 PrioSelect_77_i12_3_lut_4_lut_4_lut (.A(n11714), .B(n11_adj_1219), 
         .C(Z_N_378[0]), .D(n22248), .Z(n12_adj_1509)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_77_i12_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX mux_334_i5 (.BLUT(n1742[4]), .ALUT(n1194[4]), .C0(n1341), .Z(n1238[4]));
    LUT4 i17342_3_lut_4_lut (.A(n22219), .B(n22102), .C(n14_adj_1510), 
         .D(n10_adj_1268), .Z(n15_adj_1511)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17342_3_lut_4_lut.init = 16'hf1e0;
    PFUMX mux_334_i6 (.BLUT(n1742[5]), .ALUT(n1194[5]), .C0(n1341), .Z(n1238[5]));
    LUT4 i17694_4_lut (.A(n22157), .B(n22159), .C(n22158), .D(n213[5]), 
         .Z(n17734)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17694_4_lut.init = 16'haaab;
    LUT4 i8457_4_lut (.A(s_5_7), .B(n116), .C(n7_adj_476), .D(n7066), 
         .Z(n6_adj_1512)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i8457_4_lut.init = 16'h3022;
    LUT4 PrioSelect_77_i19_4_lut (.A(n17_adj_1513), .B(in_port[0]), .C(n9164), 
         .D(n12182), .Z(n399)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_77_i19_4_lut.init = 16'hcac0;
    LUT4 i17610_2_lut_rep_560_3_lut_4_lut_4_lut (.A(n11714), .B(n11778), 
         .C(n22277), .D(n10_adj_698), .Z(n22127)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i17610_2_lut_rep_560_3_lut_4_lut_4_lut.init = 16'h0001;
    LUT4 PrioSelect_157_i14_3_lut_4_lut (.A(n22234), .B(n11714), .C(Z_N_387[4]), 
         .D(n13_adj_1486), .Z(n14_adj_786)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_157_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_85_i12_3_lut_4_lut_4_lut (.A(n11714), .B(Z_N_367[2]), 
         .C(n1108[2]), .D(n22250), .Z(n12_adj_1514)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_85_i12_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_101_i12_3_lut_4_lut_4_lut (.A(n11714), .B(Z_N_367[6]), 
         .C(n1108[6]), .D(n22250), .Z(n12_adj_1503)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_101_i12_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_161_i14_3_lut_4_lut (.A(n22234), .B(n11714), .C(Z_N_387[5]), 
         .D(n13_adj_1474), .Z(n14_adj_793)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_161_i14_3_lut_4_lut.init = 16'hfd20;
    PFUMX mux_334_i7 (.BLUT(n1742[6]), .ALUT(n1194[6]), .C0(n1341), .Z(n1238[6]));
    LUT4 PrioSelect_165_i14_3_lut_4_lut (.A(n22234), .B(n11714), .C(Z_N_387[6]), 
         .D(n13_adj_1473), .Z(n14_adj_778)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_165_i14_3_lut_4_lut.init = 16'hfd20;
    PFUMX mux_334_i8 (.BLUT(n1742[7]), .ALUT(n1194[7]), .C0(n1341), .Z(n1238[7]));
    LUT4 i1_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), .C(n22222), 
         .D(n22106), .Z(clk_in_c_enable_16)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h3032;
    LUT4 PrioSelect_89_i12_3_lut_4_lut_4_lut (.A(n11714), .B(Z_N_367[3]), 
         .C(n1108[3]), .D(n22250), .Z(n12_adj_1515)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_89_i12_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_93_i12_3_lut_4_lut_4_lut (.A(n11714), .B(Z_N_367[4]), 
         .C(n1108[4]), .D(n22250), .Z(n12_adj_1516)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_93_i12_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_81_i12_3_lut_4_lut_4_lut (.A(n11714), .B(Z_N_367[1]), 
         .C(n1108[1]), .D(n22250), .Z(n12_adj_1517)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_81_i12_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_97_i12_3_lut_4_lut_4_lut (.A(n11714), .B(Z_N_367[5]), 
         .C(n1108[5]), .D(n22250), .Z(n12_adj_1507)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_97_i12_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_141_i14_3_lut_4_lut (.A(n22234), .B(n11714), .C(Z_N_387[0]), 
         .D(n10_adj_1471), .Z(n14_adj_978)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_141_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_169_i14_3_lut_4_lut (.A(n22234), .B(n11714), .C(Z_N_387[7]), 
         .D(n10_adj_1470), .Z(n14_adj_754)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_169_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 i14502_4_lut (.A(n22156), .B(n22155), .C(n22154), .D(n213[5]), 
         .Z(n17692)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14502_4_lut.init = 16'h5554;
    LUT4 PrioSelect_265_i8_4_lut (.A(n6_adj_1512), .B(n7_adj_473), .C(n151[5]), 
         .D(n145), .Z(n8_adj_617)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_265_i8_4_lut.init = 16'hcfca;
    LUT4 PrioSelect_77_i15_3_lut_4_lut_4_lut (.A(n11714), .B(n5), .C(n1108[0]), 
         .D(n22250), .Z(n15_adj_982)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam PrioSelect_77_i15_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 PrioSelect_493_i12_3_lut_4_lut (.A(n22258), .B(n7908), .C(Z_N_378[0]), 
         .D(n11_adj_689), .Z(n12_adj_1518)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_493_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_521_i12_3_lut_4_lut (.A(n22258), .B(n7908), .C(Z_N_378[7]), 
         .D(n11_adj_692), .Z(n12_adj_1519)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_521_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i2154_3_lut_4_lut (.A(n7762), .B(n8647), .C(n7_adj_481), .D(n7_adj_500), 
         .Z(n10_adj_883)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2154_3_lut_4_lut.init = 16'hf780;
    LUT4 i2170_3_lut_4_lut (.A(n7762), .B(n8647), .C(n7_c), .D(n7_adj_479), 
         .Z(n10_adj_900)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2170_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_334_i9 (.BLUT(n1742[8]), .ALUT(n1194[8]), .C0(n1341), .Z(n1238[8]));
    LUT4 i1498_3_lut_4_lut (.A(n8627), .B(n11714), .C(n7_c), .D(n7_adj_479), 
         .Z(n10_adj_1347)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1498_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_165 (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7908), .D(n22272), .Z(n346[15])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_165.init = 16'h0080;
    LUT4 i4_4_lut_adj_166 (.A(s_N_294[1]), .B(s_N_294[2]), .C(s_N_294[5]), 
         .D(s_N_294[4]), .Z(n10_adj_1133)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(227[81:100])
    defparam i4_4_lut_adj_166.init = 16'hfffe;
    LUT4 i1514_3_lut_4_lut (.A(n8627), .B(n11714), .C(n7_adj_462), .D(n7_adj_481), 
         .Z(n10_adj_1349)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1514_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2186_3_lut_4_lut (.A(n7762), .B(n8647), .C(n7_adj_462), .D(n7_adj_481), 
         .Z(n10_adj_895)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2186_3_lut_4_lut.init = 16'hf780;
    LUT4 i1530_3_lut_4_lut (.A(n8627), .B(n11714), .C(n7_adj_609), .D(n7_c), 
         .Z(n10_adj_1350)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1530_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17340_3_lut_4_lut (.A(n22219), .B(n22102), .C(n14_adj_1520), 
         .D(n10_adj_1262), .Z(n15_adj_1521)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17340_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17664_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22258), .B(n7908), .C(n22255), 
         .D(n22253), .Z(n19194)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17664_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hccc8;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_167 (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n11714), .D(n22272), .Z(n346[3])) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_167.init = 16'h0008;
    LUT4 PrioSelect_177_i12_3_lut_4_lut (.A(n22238), .B(n11714), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1522)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_177_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17557_4_lut (.A(n22114), .B(n22116), .C(n22115), .D(n213[15]), 
         .Z(n19574)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17557_4_lut.init = 16'haaab;
    LUT4 i17710_4_lut (.A(n22157), .B(n22159), .C(n22158), .D(n17692), 
         .Z(n20312)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17710_4_lut.init = 16'habaa;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_168 (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n16312), .D(n22272), .Z(n346[11])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_168.init = 16'h0080;
    LUT4 PrioSelect_181_i12_3_lut_4_lut (.A(n22238), .B(n11714), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1523)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_181_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_169 (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7762), .D(n22272), .Z(n346[7])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_169.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_170 (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7908), .D(n22272), .Z(n346[14])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_170.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_171 (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n16312), .D(n22272), .Z(n346[10])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_171.init = 16'h0080;
    LUT4 i8635_2_lut (.A(instruction[11]), .B(instruction[10]), .Z(n11714)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8635_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_172 (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7762), .D(n22272), .Z(n346[6])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_172.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_173 (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n11714), .D(n22272), .Z(n346[2])) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_173.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_174 (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7908), .D(n22272), .Z(n346[13])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_174.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_175 (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n16312), .D(n22272), .Z(n346[9])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_175.init = 16'h0080;
    LUT4 PrioSelect_185_i12_3_lut_4_lut (.A(n22238), .B(n11714), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1524)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_185_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2922_3_lut_4_lut (.A(n22259), .B(n7908), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1525)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i2922_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_334_i10 (.BLUT(n1742[9]), .ALUT(n1194[9]), .C0(n1341), .Z(n1238[9]));
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_176 (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7762), .D(n22272), .Z(n346[5])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_176.init = 16'h0080;
    LUT4 i17742_4_lut (.A(n22225), .B(n22224), .C(n22226), .D(n16622), 
         .Z(n20344)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam i17742_4_lut.init = 16'hefee;
    PFUMX mux_334_i11 (.BLUT(n1742[10]), .ALUT(n1194[10]), .C0(n1341), 
          .Z(n1238[10]));
    LUT4 i7_4_lut_adj_177 (.A(Z_N_387[0]), .B(n14_adj_1526), .C(n10_adj_716), 
         .D(Z_N_387[3]), .Z(C_N_351[0])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(429[15:76])
    defparam i7_4_lut_adj_177.init = 16'h6996;
    LUT4 i6_4_lut (.A(Z_N_387[5]), .B(Z_N_387[4]), .C(Z_N_387[6]), .D(Z_N_387[7]), 
         .Z(n14_adj_1526)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(429[15:76])
    defparam i6_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_178 (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n11714), .D(n22272), .Z(n346[1])) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_178.init = 16'h0008;
    PFUMX mux_334_i12 (.BLUT(n1742[11]), .ALUT(n1194[11]), .C0(n1341), 
          .Z(n1238[11]));
    LUT4 i9031_2_lut_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n11714), .D(n22272), .Z(n12182)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i9031_2_lut_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_179 (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7762), .D(n22272), .Z(n346[4])) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_179.init = 16'h0020;
    LUT4 PrioSelect_177_i17_3_lut_4_lut (.A(n7876), .B(n22220), .C(in_port[1]), 
         .D(n16_adj_1527), .Z(n17_adj_743)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_177_i17_3_lut_4_lut.init = 16'hfd20;
    PFUMX mux_334_i1 (.BLUT(n1742[0]), .ALUT(n1194[0]), .C0(n1341), .Z(n1238[0]));
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_180 (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n16312), .D(n22272), .Z(n346[8])) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_180.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_181 (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7908), .D(n22272), .Z(n346[12])) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_181.init = 16'h0020;
    LUT4 PrioSelect_189_i12_3_lut_4_lut (.A(n22238), .B(n11714), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1528)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_189_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut_4_lut_adj_182 (.A(clk_in_c_enable_174), .B(n16574), .C(n22261), 
         .D(n16375), .Z(clk_in_c_enable_94)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (C (D))) */ ;
    defparam i1_4_lut_4_lut_adj_182.init = 16'hf200;
    LUT4 i1_4_lut_4_lut_adj_183 (.A(clk_in_c_enable_174), .B(n22261), .C(n22221), 
         .D(n7762), .Z(n16378)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_adj_183.init = 16'hce00;
    LUT4 i13432_2_lut_rep_638_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n22260), 
         .C(n11916), .D(n22271), .Z(n22205)) /* synthesis lut_function=((B (C (D)))+!A) */ ;
    defparam i13432_2_lut_rep_638_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_184 (.A(clk_in_c_enable_174), .B(n22261), 
         .C(n22281), .D(n22221), .Z(clk_in_c_enable_106)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_184.init = 16'hc0e0;
    PFUMX i11646 (.BLUT(n16239), .ALUT(n16123), .C0(C), .Z(n14802));
    LUT4 PrioSelect_517_i13_3_lut_4_lut (.A(n22259), .B(n7908), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1529)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_517_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_193_i12_3_lut_4_lut (.A(n22238), .B(n11714), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1495)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_193_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_513_i13_3_lut_4_lut (.A(n22259), .B(n7908), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1530)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_513_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_509_i13_3_lut_4_lut (.A(n22259), .B(n7908), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1531)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_509_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_505_i13_3_lut_4_lut (.A(n22259), .B(n7908), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1532)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_505_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_181_i17_3_lut_4_lut (.A(n7876), .B(n22220), .C(in_port[2]), 
         .D(n16_adj_1533), .Z(n17_adj_724)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_181_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_197_i12_3_lut_4_lut (.A(n22238), .B(n11714), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1493)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_197_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_501_i13_3_lut_4_lut (.A(n22259), .B(n7908), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1534)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_501_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_185_i17_3_lut_4_lut (.A(n7876), .B(n22220), .C(in_port[3]), 
         .D(n16_adj_1535), .Z(n17_adj_691)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_185_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5_4_lut_adj_185 (.A(n16518), .B(n4_adj_1536), .C(n16520), .D(n2322), 
         .Z(n2323)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i5_4_lut_adj_185.init = 16'h0100;
    LUT4 i13357_4_lut (.A(n2319), .B(n2313), .C(n2320), .D(n2314), .Z(n16518)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i13357_4_lut.init = 16'h7bde;
    LUT4 equal_1008_i4_2_lut (.A(n2317), .B(n2318), .Z(n4_adj_1536)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(178[8] 398[4])
    defparam equal_1008_i4_2_lut.init = 16'h6666;
    LUT4 i13359_4_lut (.A(n2315), .B(n2311), .C(n2316), .D(n2312), .Z(n16520)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i13359_4_lut.init = 16'h7bde;
    LUT4 i7428_3_lut (.A(C_N_336[0]), .B(out_port_7__N_217[0]), .C(instruction[3]), 
         .Z(n103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i7428_3_lut.init = 16'hcaca;
    PFUMX PrioSelect_573_i16 (.BLUT(n11_adj_1537), .ALUT(n12_adj_1538), 
          .C0(n19547), .Z(n16_adj_1114)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_173_i15_3_lut_4_lut (.A(n22238), .B(n11714), .C(n1108[0]), 
         .D(n5_adj_1159), .Z(n15_adj_1162)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_173_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_201_i15_3_lut_4_lut (.A(n22238), .B(n11714), .C(n1108[7]), 
         .D(n9_adj_820), .Z(n15_adj_670)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_201_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_189_i17_3_lut_4_lut (.A(n7876), .B(n22220), .C(in_port[4]), 
         .D(n16_adj_1539), .Z(n17_adj_684)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_189_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_497_i13_3_lut_4_lut (.A(n22259), .B(n7908), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1540)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_497_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_193_i17_3_lut_4_lut (.A(n7876), .B(n22220), .C(in_port[5]), 
         .D(n16_adj_1496), .Z(n17_adj_680)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_193_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_197_i17_3_lut_4_lut (.A(n7876), .B(n22220), .C(in_port[6]), 
         .D(n16_adj_1494), .Z(n17_adj_677)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_197_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_521_i10_3_lut_4_lut (.A(n22259), .B(n7908), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1541)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_521_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i17558_4_lut (.A(n22116), .B(n22115), .C(n22108), .D(n19556), 
         .Z(n20160)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17558_4_lut.init = 16'hefee;
    LUT4 i1_2_lut_rep_669_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n16487), .D(n8_adj_708), .Z(n22236)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_669_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i8909_2_lut_rep_679_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n16487), .D(n8_adj_708), .Z(n22246)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i8909_2_lut_rep_679_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i16386_4_lut (.A(n22112), .B(n22113), .C(n213[15]), .D(n21255), 
         .Z(n19556)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i16386_4_lut.init = 16'h1011;
    LUT4 i2202_3_lut_4_lut (.A(n7762), .B(n8647), .C(n7_adj_609), .D(n7_c), 
         .Z(n10_adj_887)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2202_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_570_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n11714), .D(n22273), .Z(n22137)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_570_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 PrioSelect_497_i14_3_lut_4_lut (.A(n22257), .B(n7908), .C(Z_N_387[1]), 
         .D(n13_adj_1540), .Z(n14_adj_1506)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_497_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_569_i16 (.BLUT(n11_adj_1542), .ALUT(n12_adj_1543), 
          .C0(n19547), .Z(n16_adj_1112)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_153_i17_3_lut_4_lut (.A(n16392), .B(n22220), .C(in_port[3]), 
         .D(n16_adj_1544), .Z(n17_adj_816)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_153_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_501_i14_3_lut_4_lut (.A(n22257), .B(n7908), .C(Z_N_387[2]), 
         .D(n13_adj_1534), .Z(n14_adj_528)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_501_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_201_i10_3_lut_4_lut (.A(n22239), .B(n11714), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1545)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_201_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_161_i17_3_lut_4_lut (.A(n16392), .B(n22220), .C(in_port[5]), 
         .D(n16_adj_1499), .Z(n17_adj_811)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_161_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_505_i14_3_lut_4_lut (.A(n22257), .B(n7908), .C(Z_N_387[3]), 
         .D(n13_adj_1532), .Z(n14_adj_494)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_505_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_157_i17_3_lut_4_lut (.A(n16392), .B(n22220), .C(in_port[4]), 
         .D(n16_adj_1546), .Z(n17_adj_813)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_157_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_149_i17_3_lut_4_lut (.A(n16392), .B(n22220), .C(in_port[2]), 
         .D(n16_adj_1547), .Z(n17_adj_825)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_149_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17582_4_lut (.A(n22116), .B(n22115), .C(n22108), .D(n19403), 
         .Z(n20184)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17582_4_lut.init = 16'hefee;
    LUT4 i16233_4_lut (.A(n22112), .B(n22113), .C(n213[15]), .D(n19394), 
         .Z(n19403)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i16233_4_lut.init = 16'h1011;
    LUT4 n2083_bdd_4_lut_17832 (.A(n22109), .B(n2085), .C(n7762), .D(n11778), 
         .Z(n21001)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;
    defparam n2083_bdd_4_lut_17832.init = 16'hff1f;
    LUT4 PrioSelect_509_i14_3_lut_4_lut (.A(n22257), .B(n7908), .C(Z_N_387[4]), 
         .D(n13_adj_1531), .Z(n14_adj_1520)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_509_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i1802_3_lut_4_lut (.A(n22239), .B(n11714), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1548)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i1802_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_513_i14_3_lut_4_lut (.A(n22257), .B(n7908), .C(Z_N_387[5]), 
         .D(n13_adj_1530), .Z(n14_adj_1510)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_513_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_329_i8_4_lut (.A(n6_adj_1464), .B(n7_adj_473), .C(n151[7]), 
         .D(n142), .Z(n8_adj_577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_329_i8_4_lut.init = 16'hcfca;
    LUT4 PrioSelect_517_i14_3_lut_4_lut (.A(n22257), .B(n7908), .C(Z_N_387[6]), 
         .D(n13_adj_1529), .Z(n14_adj_1504)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_517_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_165_i17_3_lut_4_lut (.A(n16392), .B(n22220), .C(in_port[6]), 
         .D(n16_adj_1498), .Z(n17_adj_796)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_165_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_493_i14_3_lut_4_lut (.A(n22257), .B(n7908), .C(Z_N_387[0]), 
         .D(n10_adj_1525), .Z(n14_adj_987)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_493_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_521_i14_3_lut_4_lut (.A(n22257), .B(n7908), .C(Z_N_387[7]), 
         .D(n10_adj_1541), .Z(n14_adj_1549)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_521_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_145_i17_3_lut_4_lut (.A(n16392), .B(n22220), .C(in_port[1]), 
         .D(n16_adj_1550), .Z(n17_adj_829)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_145_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_543_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7908), .D(n22273), .Z(n22110)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_543_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_686_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n16487), .D(n8_adj_708), .Z(n22253)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_686_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i17587_4_lut (.A(n22122), .B(n22121), .C(n22107), .D(n19372), 
         .Z(n20189)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17587_4_lut.init = 16'hefee;
    LUT4 PrioSelect_113_i17_3_lut_4_lut (.A(n7726), .B(n22220), .C(in_port[1]), 
         .D(n16_adj_1551), .Z(n17_adj_875)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_113_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 i16202_4_lut (.A(n22110), .B(n22111), .C(n213[14]), .D(n21226), 
         .Z(n19372)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i16202_4_lut.init = 16'h1011;
    LUT4 PrioSelect_117_i17_3_lut_4_lut (.A(n7726), .B(n22220), .C(in_port[2]), 
         .D(n16_adj_1552), .Z(n17_adj_870)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_117_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2218_3_lut_4_lut (.A(n7762), .B(n8647), .C(n7_adj_476), .D(n7_adj_462), 
         .Z(n10_adj_898)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2218_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_197_i13_3_lut_4_lut (.A(n22239), .B(n11714), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1553)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_197_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_121_i17_3_lut_4_lut (.A(n7726), .B(n22220), .C(in_port[3]), 
         .D(n16_adj_1554), .Z(n17_adj_865)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_121_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_193_i13_3_lut_4_lut (.A(n22239), .B(n11714), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1555)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_193_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_125_i17_3_lut_4_lut (.A(n7726), .B(n22220), .C(in_port[4]), 
         .D(n16_adj_1556), .Z(n17_adj_862)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_125_i17_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_565_i16 (.BLUT(n11_adj_1557), .ALUT(n12_adj_1558), 
          .C0(n19547), .Z(n16_adj_1108)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1546_3_lut_4_lut (.A(n8627), .B(n11714), .C(n7_adj_476), .D(n7_adj_462), 
         .Z(n10_adj_1351)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i1546_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17649_4_lut (.A(n22122), .B(n22121), .C(n22107), .D(n19219), 
         .Z(n20251)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17649_4_lut.init = 16'hefee;
    LUT4 i16049_4_lut (.A(n22110), .B(n22111), .C(n213[14]), .D(n19210), 
         .Z(n19219)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i16049_4_lut.init = 16'h1011;
    PFUMX PrioSelect_561_i16 (.BLUT(n11_adj_1559), .ALUT(n12_adj_1560), 
          .C0(n19547), .Z(n16_adj_1103)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_189_i13_3_lut_4_lut (.A(n22239), .B(n11714), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1561)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_189_i13_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_21_9 (.A0(address[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(address[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14268), .COUT(n14269), .S0(n18[7]), .S1(n18[8]));   // f:/home/mini-mcu/step_fpga/mcu.v(217[27:35])
    defparam add_21_9.INIT0 = 16'h5aaa;
    defparam add_21_9.INIT1 = 16'h5aaa;
    defparam add_21_9.INJECT1_0 = "NO";
    defparam add_21_9.INJECT1_1 = "NO";
    LUT4 PrioSelect_129_i17_3_lut_4_lut (.A(n7726), .B(n22220), .C(in_port[5]), 
         .D(n16_adj_1501), .Z(n17_adj_854)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_129_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_185_i13_3_lut_4_lut (.A(n22239), .B(n11714), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1562)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_185_i13_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_541_i16 (.BLUT(n11_adj_1563), .ALUT(n12_adj_1168), 
          .C0(n19363), .Z(n16_adj_1305)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_133_i17_3_lut_4_lut (.A(n7726), .B(n22220), .C(in_port[6]), 
         .D(n16_adj_1500), .Z(n17_adj_851)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam PrioSelect_133_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2234_3_lut_4_lut (.A(n7762), .B(n8647), .C(n7_adj_473), .D(n7_adj_609), 
         .Z(n10_adj_878)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i2234_3_lut_4_lut.init = 16'hf780;
    LUT4 i17661_4_lut (.A(n22219), .B(n22218), .C(n22217), .D(n19188), 
         .Z(n20263)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17661_4_lut.init = 16'hefee;
    LUT4 PrioSelect_181_i13_3_lut_4_lut (.A(n22239), .B(n11714), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1564)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_181_i13_3_lut_4_lut.init = 16'hfd20;
    PFUMX PrioSelect_537_i16 (.BLUT(n11_adj_1565), .ALUT(n12_adj_1165), 
          .C0(n19363), .Z(n16_adj_1301)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i16018_4_lut (.A(n22216), .B(n22215), .C(n213[13]), .D(n21201), 
         .Z(n19188)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i16018_4_lut.init = 16'h1011;
    LUT4 PrioSelect_333_i5_3_lut_4_lut (.A(n8627), .B(n16312), .C(n14_adj_480), 
         .D(n14_adj_711), .Z(n5_adj_1155)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_333_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_177_i13_3_lut_4_lut (.A(n22239), .B(n11714), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1566)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_177_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17683_4_lut (.A(n22219), .B(n22218), .C(n22217), .D(n19035), 
         .Z(n20285)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17683_4_lut.init = 16'hefee;
    LUT4 i15865_4_lut (.A(n22216), .B(n22215), .C(n213[13]), .D(n19026), 
         .Z(n19035)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15865_4_lut.init = 16'h1011;
    PFUMX PrioSelect_533_i16 (.BLUT(n11_adj_1567), .ALUT(n12_adj_1164), 
          .C0(n19363), .Z(n16_adj_1299)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_594_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7762), .D(n22273), .Z(n22161)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_594_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_618_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n16312), .D(n22273), .Z(n22185)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_618_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_576_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n11714), .D(n22273), .Z(n22143)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_576_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_545_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7908), .D(n22273), .Z(n22112)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_545_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX PrioSelect_529_i16 (.BLUT(n11_adj_1568), .ALUT(n12_adj_1158), 
          .C0(n19363), .Z(n16_adj_1297)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i11184_2_lut (.A(C), .B(instruction[0]), .Z(n2055[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i11184_2_lut.init = 16'h6666;
    LUT4 PrioSelect_177_i14_3_lut_4_lut (.A(n22240), .B(n11714), .C(Z_N_387[1]), 
         .D(n13_adj_1566), .Z(n14_adj_803)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_177_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_181_i14_3_lut_4_lut (.A(n22240), .B(n11714), .C(Z_N_387[2]), 
         .D(n13_adj_1564), .Z(n14_adj_817)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_181_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_adj_186 (.A(instruction[15]), .B(instruction[13]), .Z(n4_adj_1040)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_186.init = 16'hbbbb;
    LUT4 PrioSelect_185_i14_3_lut_4_lut (.A(n22240), .B(n11714), .C(Z_N_387[3]), 
         .D(n13_adj_1562), .Z(n14_adj_807)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_185_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1307_i3_4_lut_4_lut_then_4_lut (.A(st_zc[0]), .B(st_zc[1]), 
         .C(clk_in_c_enable_109), .D(st_zc[2]), .Z(n22315)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B+((D)+!C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(206[26:38])
    defparam mux_1307_i3_4_lut_4_lut_then_4_lut.init = 16'hf7ef;
    PFUMX PrioSelect_509_i16 (.BLUT(n11_adj_685), .ALUT(n12_adj_580), .C0(n19179), 
          .Z(n16_adj_1235)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 mux_1307_i3_4_lut_4_lut_else_4_lut (.A(st_zc[0]), .B(st_zc[1]), 
         .C(clk_in_c_enable_109), .D(st_zc[2]), .Z(n22314)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B+((D)+!C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(206[26:38])
    defparam mux_1307_i3_4_lut_4_lut_else_4_lut.init = 16'h0810;
    LUT4 PrioSelect_189_i14_3_lut_4_lut (.A(n22240), .B(n11714), .C(Z_N_387[4]), 
         .D(n13_adj_1561), .Z(n14_adj_805)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_189_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 PrioSelect_193_i14_3_lut_4_lut (.A(n22240), .B(n11714), .C(Z_N_387[5]), 
         .D(n13_adj_1555), .Z(n14_adj_809)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_193_i14_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_21_7 (.A0(address[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(address[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14267), .COUT(n14268), .S0(n18[5]), .S1(n18[6]));   // f:/home/mini-mcu/step_fpga/mcu.v(217[27:35])
    defparam add_21_7.INIT0 = 16'h5aaa;
    defparam add_21_7.INIT1 = 16'h5aaa;
    defparam add_21_7.INJECT1_0 = "NO";
    defparam add_21_7.INJECT1_1 = "NO";
    PFUMX PrioSelect_505_i16 (.BLUT(n11_adj_682), .ALUT(n12_adj_563), .C0(n19179), 
          .Z(n16_adj_1233)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17530_2_lut_3_lut_4_lut (.A(n11714), .B(n22266), .C(n20131), 
         .D(n7876), .Z(n17337)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17530_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i1_2_lut_rep_600_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7762), .D(n22273), .Z(n22167)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_600_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX PrioSelect_501_i16 (.BLUT(n11_adj_678), .ALUT(n12_adj_542), .C0(n19179), 
          .Z(n16_adj_1229)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_197_i14_3_lut_4_lut (.A(n22240), .B(n11714), .C(Z_N_387[6]), 
         .D(n13_adj_1553), .Z(n14_adj_801)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_197_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 n2083_bdd_4_lut_17835 (.A(n22109), .B(n2085), .C(n7762), .D(n7726), 
         .Z(n21018)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam n2083_bdd_4_lut_17835.init = 16'h1fff;
    LUT4 PrioSelect_525_i12_3_lut_4_lut (.A(n22231), .B(n7908), .C(Z_N_378[0]), 
         .D(n11_adj_1569), .Z(n12_adj_1570)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_525_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_173_i14_3_lut_4_lut (.A(n22240), .B(n11714), .C(Z_N_387[0]), 
         .D(n10_adj_1548), .Z(n14_adj_1161)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_173_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_624_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n16312), .D(n22273), .Z(n22191)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_624_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i9039_2_lut_rep_557_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n11714), .D(n22273), .Z(n22124)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i9039_2_lut_rep_557_3_lut_4_lut_4_lut.init = 16'hfffd;
    PFUMX PrioSelect_497_i16 (.BLUT(n11_adj_681), .ALUT(n12_adj_527), .C0(n19179), 
          .Z(n16_adj_1228)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_201_i14_3_lut_4_lut (.A(n22240), .B(n11714), .C(Z_N_387[7]), 
         .D(n10_adj_1545), .Z(n14_adj_669)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_201_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_606_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n16312), .D(n22273), .Z(n22173)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_606_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 PrioSelect_553_i12_3_lut_4_lut (.A(n22231), .B(n7908), .C(Z_N_378[7]), 
         .D(n11_adj_1571), .Z(n12_adj_1572)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_553_i12_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_477_i16 (.BLUT(n11_adj_1407), .ALUT(n12_adj_1438), 
          .C0(n18995), .Z(n16_adj_1423)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17690_4_lut (.A(n22213), .B(n22212), .C(n22210), .D(n19004), 
         .Z(n20292)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17690_4_lut.init = 16'hefee;
    LUT4 i1_2_lut_rep_582_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7762), .D(n22273), .Z(n22149)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_582_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_641_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7908), .D(n22273), .Z(n22208)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_641_3_lut_4_lut_4_lut.init = 16'h0020;
    PFUMX PrioSelect_473_i16 (.BLUT(n11_adj_1406), .ALUT(n12_adj_1435), 
          .C0(n18995), .Z(n16_adj_1422)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_564_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n11714), .D(n22273), .Z(n22131)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_564_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i15834_4_lut (.A(n22208), .B(n22207), .C(n213[12]), .D(n21170), 
         .Z(n19004)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15834_4_lut.init = 16'h1011;
    LUT4 i17598_2_lut_3_lut_4_lut (.A(n11714), .B(n22266), .C(n20199), 
         .D(n16392), .Z(n17153)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17598_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i17716_2_lut_3_lut_4_lut (.A(n11714), .B(n22266), .C(n20317), 
         .D(n7726), .Z(n16969)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17716_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i1_2_lut_rep_588_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7762), .D(n22273), .Z(n22155)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_588_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 PrioSelect_213_i11_3_lut_4_lut (.A(n22245), .B(n7762), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1573)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_213_i11_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_469_i16 (.BLUT(n11_adj_1404), .ALUT(n12_adj_1434), 
          .C0(n18995), .Z(n16_adj_1421)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_612_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n16312), .D(n22273), .Z(n22179)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_612_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i17719_4_lut (.A(n22213), .B(n22212), .C(n22210), .D(n18851), 
         .Z(n20321)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17719_4_lut.init = 16'hefee;
    LUT4 i1_2_lut_rep_649_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7908), .D(n22273), .Z(n22216)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_649_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX PrioSelect_465_i16 (.BLUT(n11_adj_1405), .ALUT(n12_adj_1433), 
          .C0(n18995), .Z(n16_adj_1419)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_663_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n16487), .D(n8_adj_708), .Z(n22230)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_663_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_662_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n10_adj_586), .D(n8_adj_708), .Z(n22229)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_662_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i8846_2_lut_rep_700_3_lut_3_lut_4_lut (.A(clk_in_c_enable_174), .B(instruction[15]), 
         .C(n9_adj_707), .D(n8_adj_695), .Z(n22267)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i8846_2_lut_rep_700_3_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i15681_4_lut (.A(n22208), .B(n22207), .C(n213[12]), .D(n18842), 
         .Z(n18851)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15681_4_lut.init = 16'h1011;
    PFUMX PrioSelect_445_i16 (.BLUT(n11_adj_1263), .ALUT(n12_adj_1277), 
          .C0(n18811), .Z(n16_adj_1314)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_544_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7908), .D(n22274), .Z(n22111)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_544_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i13434_2_lut_rep_539_4_lut (.A(n22271), .B(n11916), .C(n22260), 
         .D(n11714), .Z(n22106)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i13434_2_lut_rep_539_4_lut.init = 16'hff80;
    LUT4 PrioSelect_209_i11_3_lut_4_lut (.A(n22245), .B(n7762), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1574)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_209_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_668_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n10_adj_586), .D(n8_adj_708), .Z(n22235)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_668_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 n2083_bdd_4_lut_17847 (.A(n22109), .B(n2085), .C(n7762), .D(n7876), 
         .Z(n21062)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam n2083_bdd_4_lut_17847.init = 16'h1fff;
    PFUMX PrioSelect_441_i16 (.BLUT(n11_adj_1261), .ALUT(n12_adj_1283), 
          .C0(n18811), .Z(n16_adj_1313)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_631_4_lut (.A(n22271), .B(n11916), .C(n22260), .D(n22280), 
         .Z(n22198)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(D))) */ ;
    defparam i1_2_lut_rep_631_4_lut.init = 16'h7f00;
    LUT4 PrioSelect_217_i11_3_lut_4_lut (.A(n22245), .B(n7762), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1575)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_217_i11_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_437_i16 (.BLUT(n11_adj_1258), .ALUT(n12_adj_1281), 
          .C0(n18811), .Z(n16_adj_1312)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i8901_2_lut_rep_678_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n10_adj_586), .D(n8_adj_708), .Z(n22245)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i8901_2_lut_rep_678_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_rep_569_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n11714), .D(n22274), .Z(n22136)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_569_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_593_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7762), .D(n22274), .Z(n22160)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_593_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_617_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n16312), .D(n22274), .Z(n22184)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_617_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_546_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7908), .D(n22274), .Z(n22113)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_546_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 PrioSelect_393_i8_4_lut (.A(n6_adj_1446), .B(n14_adj_711), .C(n16326), 
         .D(n16346), .Z(n8_adj_543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_393_i8_4_lut.init = 16'hcfca;
    LUT4 i1_2_lut_rep_688_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n10_adj_586), .D(n8_adj_708), .Z(n22255)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_688_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_575_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n11714), .D(n22274), .Z(n22142)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_575_3_lut_4_lut_4_lut.init = 16'h0008;
    PFUMX PrioSelect_433_i16 (.BLUT(n11_adj_1259), .ALUT(n12_adj_1280), 
          .C0(n18811), .Z(n16_adj_1311)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_599_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7762), .D(n22274), .Z(n22166)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_599_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 PrioSelect_221_i11_3_lut_4_lut (.A(n22245), .B(n7762), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1576)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_221_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_623_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n16312), .D(n22274), .Z(n22190)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_623_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX PrioSelect_413_i16 (.BLUT(n11_adj_1223), .ALUT(n12_adj_1245), 
          .C0(n18627), .Z(n16_adj_1321)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17722_4_lut (.A(n22195), .B(n22194), .C(n22192), .D(n18820), 
         .Z(n20324)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17722_4_lut.init = 16'hefee;
    LUT4 i15650_4_lut (.A(n22191), .B(n22190), .C(n213[11]), .D(n21132), 
         .Z(n18820)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15650_4_lut.init = 16'h1011;
    LUT4 PrioSelect_557_i12_3_lut_4_lut (.A(n22237), .B(n7908), .C(Z_N_378[0]), 
         .D(n11_adj_1577), .Z(n12_adj_1578)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_557_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i17625_2_lut_rep_556_3_lut_4_lut_4_lut_4_lut (.A(clk_in_c_enable_174), 
         .B(n22274), .C(n11778), .D(n11714), .Z(n22123)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i17625_2_lut_rep_556_3_lut_4_lut_4_lut_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_605_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n16312), .D(n22274), .Z(n22172)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_605_3_lut_4_lut_4_lut.init = 16'h0020;
    PFUMX PrioSelect_409_i16 (.BLUT(n11_adj_1222), .ALUT(n12_adj_1244), 
          .C0(n18627), .Z(n16_adj_1320)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17756_4_lut (.A(n22195), .B(n22194), .C(n22192), .D(n18667), 
         .Z(n20358)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17756_4_lut.init = 16'hefee;
    LUT4 i15497_4_lut (.A(n22191), .B(n22190), .C(n213[11]), .D(n18658), 
         .Z(n18667)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15497_4_lut.init = 16'h1011;
    PFUMX PrioSelect_405_i16 (.BLUT(n11_adj_1220), .ALUT(n12_adj_1243), 
          .C0(n18627), .Z(n16_adj_1319)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_225_i11_3_lut_4_lut (.A(n22245), .B(n7762), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1489)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_225_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_640_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7908), .D(n22274), .Z(n22207)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_640_3_lut_4_lut_4_lut.init = 16'h0020;
    PFUMX PrioSelect_401_i16 (.BLUT(n11_adj_1221), .ALUT(n12_adj_1240), 
          .C0(n18627), .Z(n16_adj_1318)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_581_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7762), .D(n22274), .Z(n22148)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_581_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_563_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n11714), .D(n22274), .Z(n22130)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_563_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 C_N_340_7__I_0_587_i15_2_lut_rep_656 (.A(C_N_336[0]), .B(C_N_342[7]), 
         .Z(n22223)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam C_N_340_7__I_0_587_i15_2_lut_rep_656.init = 16'h6666;
    PFUMX PrioSelect_381_i16 (.BLUT(n11_adj_1189), .ALUT(n12_adj_1203), 
          .C0(n18363), .Z(n16_adj_1327)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_585_i12_3_lut_4_lut (.A(n22237), .B(n7908), .C(Z_N_378[7]), 
         .D(n11_adj_1579), .Z(n12_adj_1580)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_585_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 C_N_340_7__I_0_587_i12_3_lut_3_lut (.A(C_N_336[0]), .B(C_N_342[7]), 
         .C(n10_adj_1581), .Z(n12_adj_1582)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam C_N_340_7__I_0_587_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 PrioSelect_229_i11_3_lut_4_lut (.A(n22245), .B(n7762), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1484)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_229_i11_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_377_i16 (.BLUT(n11_adj_1188), .ALUT(n12_adj_1202), 
          .C0(n18363), .Z(n16_adj_1326)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17759_4_lut (.A(n22189), .B(n22188), .C(n22186), .D(n18636), 
         .Z(n20361)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17759_4_lut.init = 16'hefee;
    LUT4 i15466_4_lut (.A(n22185), .B(n22184), .C(n213[10]), .D(n21115), 
         .Z(n18636)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15466_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_rep_587_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7762), .D(n22274), .Z(n22154)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_587_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX PrioSelect_373_i16 (.BLUT(n11_adj_1179), .ALUT(n12_adj_1201), 
          .C0(n18363), .Z(n16_adj_1325)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_611_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n16312), .D(n22274), .Z(n22178)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_611_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_648_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7908), .D(n22274), .Z(n22215)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_648_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_187 (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7908), .D(n22275), .Z(n213[14])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_187.init = 16'h0080;
    LUT4 i8899_2_lut_rep_682_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n10_adj_586), .D(n8_adj_849), .Z(n22249)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i8899_2_lut_rep_682_3_lut_4_lut_4_lut.init = 16'hfffd;
    PFUMX PrioSelect_369_i16 (.BLUT(n11_adj_1186), .ALUT(n12_adj_1200), 
          .C0(n18363), .Z(n16_adj_1324)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_188 (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7762), .D(n22275), .Z(n213[6])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_188.init = 16'h0080;
    LUT4 i17743_2_lut_3_lut (.A(C_N_336[0]), .B(C_N_342[7]), .C(n20344), 
         .Z(n16636)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam i17743_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i17775_4_lut (.A(n22189), .B(n22188), .C(n22186), .D(n18483), 
         .Z(n20377)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17775_4_lut.init = 16'hefee;
    LUT4 i15313_4_lut (.A(n22185), .B(n22184), .C(n213[10]), .D(n18474), 
         .Z(n18483)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15313_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_189 (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n11714), .D(n22275), .Z(n213[2])) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_189.init = 16'h0008;
    PFUMX PrioSelect_349_i16 (.BLUT(n11_adj_1139), .ALUT(n12_adj_1152), 
          .C0(n18259), .Z(n16_adj_1334)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_525_i11_3_lut_4_lut (.A(n22230), .B(n7908), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1569)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_525_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_190 (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n16312), .D(n22275), .Z(n213[10])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_190.init = 16'h0080;
    LUT4 C_N_340_7__I_0_587_i11_2_lut_rep_657 (.A(s_N_294[5]), .B(C_N_342[5]), 
         .Z(n22224)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam C_N_340_7__I_0_587_i11_2_lut_rep_657.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_191 (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7908), .D(n22275), .Z(n213[15])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_191.init = 16'h0080;
    CCU2D add_412_9 (.A0(instruction[7]), .B0(instruction[11]), .C0(n7_adj_473), 
          .D0(n14_adj_711), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14277), .S0(Z_N_378[7]), .S1(n1384));   // f:/home/mini-mcu/step_fpga/mcu.v(275[74:85])
    defparam add_412_9.INIT0 = 16'ha965;
    defparam add_412_9.INIT1 = 16'h0000;
    defparam add_412_9.INJECT1_0 = "NO";
    defparam add_412_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_192 (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n11714), .D(n22275), .Z(n213[3])) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_192.init = 16'h0008;
    PFUMX PrioSelect_345_i16 (.BLUT(n11_adj_1138), .ALUT(n12_adj_1151), 
          .C0(n18259), .Z(n16_adj_1333)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 C_N_340_7__I_0_587_i13_2_lut_rep_658 (.A(s_N_294[6]), .B(C_N_342[6]), 
         .Z(n22225)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam C_N_340_7__I_0_587_i13_2_lut_rep_658.init = 16'h6666;
    LUT4 i13463_2_lut_3_lut_4_lut (.A(s_N_294[6]), .B(C_N_342[6]), .C(C_N_342[5]), 
         .D(s_N_294[5]), .Z(n16633)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam i13463_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 C_N_340_7__I_0_587_i10_3_lut_3_lut (.A(s_N_294[6]), .B(C_N_342[6]), 
         .C(C_N_342[5]), .Z(n10_adj_1581)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam C_N_340_7__I_0_587_i10_3_lut_3_lut.init = 16'hd4d4;
    PFUMX PrioSelect_341_i16 (.BLUT(n11_adj_1136), .ALUT(n12_adj_1150), 
          .C0(n18259), .Z(n16_adj_1332)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_193 (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n16312), .D(n22275), .Z(n213[11])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_193.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_194 (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7762), .D(n22275), .Z(n213[7])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_194.init = 16'h0080;
    PFUMX PrioSelect_337_i16 (.BLUT(n11_adj_1137), .ALUT(n12_adj_1149), 
          .C0(n18259), .Z(n16_adj_1331)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17780_4_lut (.A(n22183), .B(n22182), .C(n22180), .D(n18452), 
         .Z(n20382)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17780_4_lut.init = 16'hefee;
    LUT4 PrioSelect_553_i11_3_lut_4_lut (.A(n22230), .B(n7908), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1571)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_553_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i15282_4_lut (.A(n22179), .B(n22178), .C(n213[9]), .D(n21098), 
         .Z(n18452)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15282_4_lut.init = 16'h1011;
    LUT4 i9026_2_lut_rep_559_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n11714), .D(n22275), .Z(n22126)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i9026_2_lut_rep_559_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 PrioSelect_233_i11_3_lut_4_lut (.A(n22246), .B(n7762), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1583)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_233_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_533_i11_3_lut_4_lut (.A(n22229), .B(n7908), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1567)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_533_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_317_i16 (.BLUT(n11_adj_1023), .ALUT(n12_adj_1070), 
          .C0(n18075), .Z(n16_adj_1341)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    CCU2D add_412_7 (.A0(instruction[5]), .B0(instruction[11]), .C0(n7_adj_609), 
          .D0(n14_adj_705), .A1(instruction[6]), .B1(instruction[11]), 
          .C1(n7_adj_476), .D1(n14_adj_709), .CIN(n14276), .COUT(n14277), 
          .S0(Z_N_378[5]), .S1(Z_N_378[6]));   // f:/home/mini-mcu/step_fpga/mcu.v(275[74:85])
    defparam add_412_7.INIT0 = 16'ha965;
    defparam add_412_7.INIT1 = 16'ha965;
    defparam add_412_7.INJECT1_0 = "NO";
    defparam add_412_7.INJECT1_1 = "NO";
    LUT4 C_N_340_7__I_0_587_i6_3_lut_3_lut (.A(s_N_294[3]), .B(C_N_342[3]), 
         .C(C_N_342[2]), .Z(n6_adj_1584)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam C_N_340_7__I_0_587_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_195 (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7908), .D(n22275), .Z(n213[12])) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_195.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_196 (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n16312), .D(n22275), .Z(n213[8])) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_196.init = 16'h0020;
    LUT4 i17493_4_lut (.A(n22183), .B(n22182), .C(n22180), .D(n18299), 
         .Z(n20095)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17493_4_lut.init = 16'hefee;
    LUT4 i15129_4_lut (.A(n22179), .B(n22178), .C(n213[9]), .D(n18290), 
         .Z(n18299)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15129_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_197 (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7762), .D(n22275), .Z(n213[4])) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_197.init = 16'h0020;
    PFUMX PrioSelect_313_i16 (.BLUT(n11_adj_1017), .ALUT(n12_adj_1066), 
          .C0(n18075), .Z(n16_adj_1340)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_198 (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7762), .D(n22275), .Z(n213[5])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_198.init = 16'h0080;
    LUT4 i13452_3_lut_4_lut (.A(s_N_294[3]), .B(C_N_342[3]), .C(C_N_342[2]), 
         .D(s_N_294[2]), .Z(n16622)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam i13452_3_lut_4_lut.init = 16'h9009;
    LUT4 PrioSelect_205_i11_3_lut_4_lut (.A(n22246), .B(n7762), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1585)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_205_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_529_i11_3_lut_4_lut (.A(n22229), .B(n7908), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1568)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_529_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_309_i16 (.BLUT(n11_adj_999), .ALUT(n12_adj_1065), .C0(n18075), 
          .Z(n16_adj_1339)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 C_N_340_7__I_0_587_i9_2_lut_rep_659 (.A(s_N_294[4]), .B(C_N_342[4]), 
         .Z(n22226)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam C_N_340_7__I_0_587_i9_2_lut_rep_659.init = 16'h6666;
    LUT4 C_N_340_7__I_0_587_i8_3_lut_3_lut (.A(s_N_294[4]), .B(C_N_342[4]), 
         .C(n6_adj_1584), .Z(n8_adj_1416)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam C_N_340_7__I_0_587_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_199 (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n11714), .D(n22275), .Z(n213[1])) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_199.init = 16'h0008;
    PFUMX PrioSelect_305_i16 (.BLUT(n11_adj_1014), .ALUT(n12_adj_1064), 
          .C0(n18075), .Z(n16_adj_1338)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i229_2_lut (.A(instruction[1]), .B(instruction[2]), .Z(n206)) /* synthesis lut_function=(A (B)) */ ;
    defparam i229_2_lut.init = 16'h8888;
    LUT4 PrioSelect_537_i11_3_lut_4_lut (.A(n22229), .B(n7908), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1565)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_537_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_200 (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n16312), .D(n22275), .Z(n213[9])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_200.init = 16'h0080;
    LUT4 PrioSelect_541_i11_3_lut_4_lut (.A(n22229), .B(n7908), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1563)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_541_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_285_i16 (.BLUT(n11_adj_764), .ALUT(n12_adj_908), .C0(n17891), 
          .Z(n16_adj_1355)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_545_i11_3_lut_4_lut (.A(n22229), .B(n7908), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1445)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_545_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_201 (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7908), .D(n22275), .Z(n213[13])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_201.init = 16'h0080;
    LUT4 PrioSelect_549_i11_3_lut_4_lut (.A(n22229), .B(n7908), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1443)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_549_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_281_i16 (.BLUT(n11_adj_763), .ALUT(n12_adj_909), .C0(n17891), 
          .Z(n16_adj_1354)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17526_4_lut (.A(n22177), .B(n22176), .C(n22174), .D(n18268), 
         .Z(n20128)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17526_4_lut.init = 16'hefee;
    LUT4 i17590_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22229), .B(n7908), .C(n22231), 
         .D(n22230), .Z(n19378)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam i17590_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hccc8;
    PFUMX PrioSelect_277_i16 (.BLUT(n11_adj_746), .ALUT(n12_adj_918), .C0(n17891), 
          .Z(n16_adj_1348)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i15098_4_lut (.A(n22173), .B(n22172), .C(n213[8]), .D(n21081), 
         .Z(n18268)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i15098_4_lut.init = 16'h1011;
    LUT4 i17755_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22248), .B(n7762), .C(n22245), 
         .D(n22246), .Z(n17538)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17755_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h4ccc;
    PFUMX PrioSelect_273_i16 (.BLUT(n11_adj_753), .ALUT(n12_adj_919), .C0(n17891), 
          .Z(n16_adj_1352)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17553_4_lut (.A(n22177), .B(n22176), .C(n22174), .D(n18115), 
         .Z(n20155)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17553_4_lut.init = 16'hefee;
    LUT4 i14945_4_lut (.A(n22173), .B(n22172), .C(n213[8]), .D(n18106), 
         .Z(n18115)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14945_4_lut.init = 16'h1011;
    LUT4 PrioSelect_233_i12_3_lut_4_lut (.A(n22248), .B(n7762), .C(Z_N_378[7]), 
         .D(n11_adj_1583), .Z(n12_adj_1586)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_233_i12_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_253_i16 (.BLUT(n11_adj_1587), .ALUT(n12_adj_1588), 
          .C0(n17707), .Z(n16_adj_1363)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i13438_2_lut_rep_653_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), 
         .B(n8050), .C(n11714), .D(n10_adj_698), .Z(n22220)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i13438_2_lut_rep_653_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 PrioSelect_557_i11_3_lut_4_lut (.A(n22236), .B(n7908), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1577)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_557_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_205_i12_3_lut_4_lut (.A(n22248), .B(n7762), .C(Z_N_378[0]), 
         .D(n11_adj_1585), .Z(n12_adj_1589)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_205_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17565_4_lut (.A(n22171), .B(n22170), .C(n22168), .D(n18084), 
         .Z(n20167)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17565_4_lut.init = 16'hefee;
    LUT4 i1_2_lut_rep_674_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n8050), 
         .C(n22281), .D(n10_adj_698), .Z(n22241)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_674_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_675_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n8050), 
         .C(n16312), .D(n10_adj_698), .Z(n22242)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_675_3_lut_4_lut_4_lut.init = 16'h0020;
    PFUMX PrioSelect_249_i16 (.BLUT(n11_adj_1590), .ALUT(n12_adj_1591), 
          .C0(n17707), .Z(n16_adj_1362)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i14914_4_lut (.A(n22167), .B(n22166), .C(n213[7]), .D(n21062), 
         .Z(n18084)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14914_4_lut.init = 16'h1011;
    LUT4 PrioSelect_105_i19_4_lut (.A(n17_adj_1592), .B(in_port[7]), .C(n9164), 
         .D(n12182), .Z(n427)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_105_i19_4_lut.init = 16'hcac0;
    LUT4 PrioSelect_585_i11_3_lut_4_lut (.A(n22236), .B(n7908), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1579)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_585_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i17601_4_lut (.A(n22171), .B(n22170), .C(n22168), .D(n17931), 
         .Z(n20203)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17601_4_lut.init = 16'hefee;
    LUT4 i14761_4_lut (.A(n22167), .B(n22166), .C(n213[7]), .D(n17922), 
         .Z(n17931)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14761_4_lut.init = 16'h1011;
    LUT4 PrioSelect_109_i19_4_lut (.A(n17_adj_1593), .B(in_port[0]), .C(n22105), 
         .D(n346[1]), .Z(n431)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_109_i19_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_rep_677_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n8050), 
         .C(n7762), .D(n10_adj_698), .Z(n22244)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_677_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_680_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n8050), 
         .C(n7908), .D(n10_adj_698), .Z(n22247)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_680_3_lut_4_lut_4_lut.init = 16'h0020;
    PFUMX PrioSelect_245_i16 (.BLUT(n11_adj_1594), .ALUT(n12_adj_1595), 
          .C0(n17707), .Z(n16_adj_1359)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_689_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n8050), 
         .C(n16375), .D(n10_adj_698), .Z(n22256)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_689_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 PrioSelect_209_i12_3_lut_4_lut (.A(n22250), .B(n7762), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1596)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_209_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_565_i11_3_lut_4_lut (.A(n22235), .B(n7908), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1557)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_565_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_241_i16 (.BLUT(n11_adj_1597), .ALUT(n12_adj_1598), 
          .C0(n17707), .Z(n16_adj_1358)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_561_i11_3_lut_4_lut (.A(n22235), .B(n7908), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1559)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_561_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_569_i11_3_lut_4_lut (.A(n22235), .B(n7908), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1542)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_569_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i17629_4_lut (.A(n22165), .B(n22164), .C(n22162), .D(n17900), 
         .Z(n20231)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17629_4_lut.init = 16'hefee;
    LUT4 PrioSelect_213_i12_3_lut_4_lut (.A(n22250), .B(n7762), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1599)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_213_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i14730_4_lut (.A(n22161), .B(n22160), .C(n213[6]), .D(n21035), 
         .Z(n17900)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14730_4_lut.init = 16'h1011;
    PFUMX PrioSelect_221_i16 (.BLUT(n11_adj_1576), .ALUT(n12_adj_1600), 
          .C0(n17523), .Z(n16_adj_1401)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_573_i11_3_lut_4_lut (.A(n22235), .B(n7908), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1537)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_573_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_217_i12_3_lut_4_lut (.A(n22250), .B(n7762), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1601)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_217_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_221_i12_3_lut_4_lut (.A(n22250), .B(n7762), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1600)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_221_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_225_i12_3_lut_4_lut (.A(n22250), .B(n7762), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1490)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_225_i12_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_217_i16 (.BLUT(n11_adj_1575), .ALUT(n12_adj_1601), 
          .C0(n17523), .Z(n16_adj_1400)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17685_4_lut (.A(n22165), .B(n22164), .C(n22162), .D(n17747), 
         .Z(n20287)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17685_4_lut.init = 16'hefee;
    LUT4 i14577_4_lut (.A(n22161), .B(n22160), .C(n213[6]), .D(n17738), 
         .Z(n17747)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14577_4_lut.init = 16'h1011;
    PFUMX i18417 (.BLUT(n22326), .ALUT(n22327), .C0(instruction[12]), 
          .Z(n22328));
    LUT4 i1_2_lut_rep_665_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n10_adj_698), 
         .C(n16392), .D(n8_adj_695), .Z(n22232)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_665_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 PrioSelect_229_i12_3_lut_4_lut (.A(n22250), .B(n7762), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1485)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_229_i12_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_213_i16 (.BLUT(n11_adj_1573), .ALUT(n12_adj_1599), 
          .C0(n17523), .Z(n16_adj_1392)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_671_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n10_adj_698), 
         .C(n7876), .D(n8_adj_695), .Z(n22238)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_671_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 n2083_bdd_4_lut_17838 (.A(n22109), .B(n2085), .C(n7762), .D(n16392), 
         .Z(n21035)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam n2083_bdd_4_lut_17838.init = 16'h1fff;
    LUT4 i8895_2_lut_rep_683_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n10_adj_698), 
         .C(n11778), .D(n8_adj_695), .Z(n22250)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i8895_2_lut_rep_683_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_rep_687_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n10_adj_698), 
         .C(n7726), .D(n8_adj_695), .Z(n22254)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_687_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_667_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n10_adj_586), 
         .C(n16392), .D(n8_adj_695), .Z(n22234)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_667_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i6951_1_lut_rep_661 (.A(out_port_7__N_217[0]), .Z(n22228)) /* synthesis lut_function=(!(A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(406[24:28])
    defparam i6951_1_lut_rep_661.init = 16'h5555;
    LUT4 C_N_340_7__I_0_587_i4_4_lut_4_lut (.A(out_port_7__N_217[0]), .B(s_N_294[1]), 
         .C(C_N_342[1]), .D(n2055[0]), .Z(n4_adj_1602)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C (D))+!B (C+(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(406[24:28])
    defparam C_N_340_7__I_0_587_i4_4_lut_4_lut.init = 16'h7130;
    LUT4 PrioSelect_577_i11_3_lut_4_lut (.A(n22235), .B(n7908), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1439)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_577_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_205_i15_3_lut_4_lut (.A(n22250), .B(n7762), .C(n1108[0]), 
         .D(n5_adj_1429), .Z(n15_adj_974)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_205_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_673_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n10_adj_586), 
         .C(n7876), .D(n8_adj_695), .Z(n22240)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_673_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 PrioSelect_581_i11_3_lut_4_lut (.A(n22235), .B(n7908), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1436)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_581_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i17561_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22235), .B(n7908), .C(n22237), 
         .D(n22236), .Z(n19562)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam i17561_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hccc8;
    LUT4 i8907_2_lut_rep_684_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n10_adj_586), 
         .C(n11778), .D(n8_adj_695), .Z(n22251)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i8907_2_lut_rep_684_3_lut_4_lut_4_lut.init = 16'hfffd;
    PFUMX PrioSelect_209_i16 (.BLUT(n11_adj_1574), .ALUT(n12_adj_1596), 
          .C0(n17523), .Z(n16_adj_1383)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_690_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n10_adj_586), 
         .C(n7726), .D(n8_adj_695), .Z(n22257)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_690_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i17042_4_lut_4_lut (.A(n22223), .B(n16633), .C(n12_adj_1582), 
         .D(n4_adj_1602), .Z(n14_adj_1417)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[80:113])
    defparam i17042_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_666_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n10_adj_863), .D(n8_adj_695), .Z(n22233)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_666_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_554_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7908), .D(n22278), .Z(n22121)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_554_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX i18085 (.BLUT(n21531), .ALUT(n21530), .C0(instruction[17]), 
          .Z(n21532));
    LUT4 i8897_2_lut_rep_685_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n10_adj_863), .D(n8_adj_695), .Z(n22252)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i8897_2_lut_rep_685_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_rep_672_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n10_adj_863), .D(n8_adj_695), .Z(n22239)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_672_3_lut_4_lut_4_lut.init = 16'h0008;
    PFUMX PrioSelect_189_i16 (.BLUT(n11_adj_664), .ALUT(n12_adj_1528), .C0(n17339), 
          .Z(n16_adj_1539)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_233_i15_3_lut_4_lut (.A(n22250), .B(n7762), .C(n1108[7]), 
         .D(n9_adj_864), .Z(n15_adj_640)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_233_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17695_4_lut (.A(n22159), .B(n22158), .C(n22156), .D(n17716), 
         .Z(n20297)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17695_4_lut.init = 16'hefee;
    LUT4 i14546_4_lut (.A(n22155), .B(n22154), .C(n213[5]), .D(n21018), 
         .Z(n17716)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14546_4_lut.init = 16'h1011;
    PFUMX PrioSelect_185_i16 (.BLUT(n11_adj_663), .ALUT(n12_adj_1524), .C0(n17339), 
          .Z(n16_adj_1535)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_573_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n11714), .D(n22278), .Z(n22140)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_573_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i17744_4_lut (.A(n22159), .B(n22158), .C(n22156), .D(n17563), 
         .Z(n20346)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17744_4_lut.init = 16'hefee;
    LUT4 i14393_4_lut (.A(n22155), .B(n22154), .C(n213[5]), .D(n17554), 
         .Z(n17563)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14393_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_rep_597_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7762), .D(n22278), .Z(n22164)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_597_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 PrioSelect_233_i10_3_lut_4_lut (.A(n22252), .B(n7762), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1603)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_233_i10_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_181_i16 (.BLUT(n11_adj_519), .ALUT(n12_adj_1523), .C0(n17339), 
          .Z(n16_adj_1533)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_621_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n16312), .D(n22278), .Z(n22188)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_621_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 PrioSelect_561_i12_3_lut_4_lut (.A(n22238), .B(n7908), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1560)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_561_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_548_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7908), .D(n22278), .Z(n22115)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_548_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX PrioSelect_177_i16 (.BLUT(n11_adj_654), .ALUT(n12_adj_1522), .C0(n17339), 
          .Z(n16_adj_1527)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1914_3_lut_4_lut (.A(n22252), .B(n7762), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1604)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i1914_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_579_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n11714), .D(n22278), .Z(n22146)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_579_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 PrioSelect_565_i12_3_lut_4_lut (.A(n22238), .B(n7908), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1558)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_565_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_229_i13_3_lut_4_lut (.A(n22252), .B(n7762), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1605)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_229_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_569_i12_3_lut_4_lut (.A(n22238), .B(n7908), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1543)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_569_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_603_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7762), .D(n22278), .Z(n22170)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_603_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_627_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n16312), .D(n22278), .Z(n22194)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_627_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_692_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n10_adj_863), .D(n8_adj_695), .Z(n22259)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_692_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i9024_2_lut_rep_561_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n11714), .D(n22278), .Z(n22128)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i9024_2_lut_rep_561_3_lut_4_lut_4_lut.init = 16'hfffd;
    PFUMX PrioSelect_157_i16 (.BLUT(n11_adj_1418), .ALUT(n12_adj_1465), 
          .C0(n17155), .Z(n16_adj_1546)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17752_4_lut (.A(n22153), .B(n22152), .C(n22150), .D(n17532), 
         .Z(n20354)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17752_4_lut.init = 16'hefee;
    LUT4 PrioSelect_573_i12_3_lut_4_lut (.A(n22238), .B(n7908), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1538)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_573_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i14362_4_lut (.A(n22149), .B(n22148), .C(n213[4]), .D(n21001), 
         .Z(n17532)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14362_4_lut.init = 16'h1011;
    LUT4 PrioSelect_225_i13_3_lut_4_lut (.A(n22252), .B(n7762), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1606)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_225_i13_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_153_i16 (.BLUT(n11_adj_1414), .ALUT(n12_adj_1468), 
          .C0(n17155), .Z(n16_adj_1544)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_221_i13_3_lut_4_lut (.A(n22252), .B(n7762), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1607)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_221_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17782_4_lut (.A(n22153), .B(n22152), .C(n22150), .D(n17379), 
         .Z(n20384)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17782_4_lut.init = 16'hefee;
    PFUMX PrioSelect_149_i16 (.BLUT(n11_adj_1412), .ALUT(n12_adj_1463), 
          .C0(n17155), .Z(n16_adj_1547)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i14209_4_lut (.A(n22149), .B(n22148), .C(n213[4]), .D(n17370), 
         .Z(n17379)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14209_4_lut.init = 16'h1011;
    LUT4 PrioSelect_217_i13_3_lut_4_lut (.A(n22252), .B(n7762), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1608)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_217_i13_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_145_i16 (.BLUT(n11_adj_1413), .ALUT(n12_adj_1467), 
          .C0(n17155), .Z(n16_adj_1550)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_213_i13_3_lut_4_lut (.A(n22252), .B(n7762), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1609)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_213_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_209_i13_3_lut_4_lut (.A(n22252), .B(n7762), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1610)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_209_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_577_i12_3_lut_4_lut (.A(n22238), .B(n7908), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1440)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_577_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_585_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7762), .D(n22278), .Z(n22152)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_585_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 PrioSelect_209_i14_3_lut_4_lut (.A(n22251), .B(n7762), .C(Z_N_387[1]), 
         .D(n13_adj_1610), .Z(n14_adj_823)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_209_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_609_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n16312), .D(n22278), .Z(n22176)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_609_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 PrioSelect_581_i12_3_lut_4_lut (.A(n22238), .B(n7908), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1437)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_581_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_213_i14_3_lut_4_lut (.A(n22251), .B(n7762), .C(Z_N_387[2]), 
         .D(n13_adj_1609), .Z(n14_adj_857)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_213_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_217_i14_3_lut_4_lut (.A(n22251), .B(n7762), .C(Z_N_387[3]), 
         .D(n13_adj_1608), .Z(n14_adj_831)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_217_i14_3_lut_4_lut.init = 16'hfb40;
    PFUMX PrioSelect_125_i16 (.BLUT(n11_adj_1285), .ALUT(n12_adj_1343), 
          .C0(n16971), .Z(n16_adj_1556)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_645_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7908), .D(n22278), .Z(n22212)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_645_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 PrioSelect_137_i19_4_lut (.A(n17_adj_1611), .B(in_port[7]), .C(n22105), 
         .D(n346[1]), .Z(n459)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_137_i19_4_lut.init = 16'hc0ca;
    LUT4 PrioSelect_221_i14_3_lut_4_lut (.A(n22251), .B(n7762), .C(Z_N_387[4]), 
         .D(n13_adj_1607), .Z(n14_adj_826)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_221_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_567_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n11714), .D(n22278), .Z(n22134)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_567_3_lut_4_lut_4_lut.init = 16'h0008;
    PFUMX PrioSelect_121_i16 (.BLUT(n11_adj_1282), .ALUT(n12_adj_1342), 
          .C0(n16971), .Z(n16_adj_1554)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_557_i15_3_lut_4_lut (.A(n22238), .B(n7908), .C(n1108[0]), 
         .D(n5_adj_1612), .Z(n15_adj_1216)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_557_i15_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_117_i16 (.BLUT(n11_adj_1276), .ALUT(n12_adj_1337), 
          .C0(n16971), .Z(n16_adj_1552)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_141_i19_4_lut (.A(n17_adj_1613), .B(in_port[0]), .C(n22104), 
         .D(n346[2]), .Z(n463)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_141_i19_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_rep_591_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7762), .D(n22278), .Z(n22158)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_591_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_615_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n16312), .D(n22278), .Z(n22182)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_615_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 PrioSelect_585_i15_3_lut_4_lut (.A(n22238), .B(n7908), .C(n1108[7]), 
         .D(n9_adj_1466), .Z(n15_adj_1614)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_585_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_651_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7908), .D(n22278), .Z(n22218)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_651_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i17475_4_lut (.A(n22147), .B(n22146), .C(n22144), .D(n17348), 
         .Z(n20077)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17475_4_lut.init = 16'hefee;
    LUT4 i14178_4_lut (.A(n22143), .B(n22142), .C(n213[3]), .D(n20976), 
         .Z(n17348)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14178_4_lut.init = 16'h1011;
    LUT4 PrioSelect_581_i13_3_lut_4_lut (.A(n22239), .B(n7908), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_1615)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_581_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i17562_4_lut (.A(n22147), .B(n22146), .C(n22144), .D(n17195), 
         .Z(n20164)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17562_4_lut.init = 16'hefee;
    LUT4 PrioSelect_225_i14_3_lut_4_lut (.A(n22251), .B(n7762), .C(Z_N_387[5]), 
         .D(n13_adj_1606), .Z(n14_adj_835)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_225_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i14025_4_lut (.A(n22143), .B(n22142), .C(n213[3]), .D(n17186), 
         .Z(n17195)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i14025_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_rep_540_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7908), .D(n22279), .Z(n22107)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_540_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX PrioSelect_113_i16 (.BLUT(n11_adj_1278), .ALUT(n12_adj_1330), 
          .C0(n16971), .Z(n16_adj_1551)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_229_i14_3_lut_4_lut (.A(n22251), .B(n7762), .C(Z_N_387[6]), 
         .D(n13_adj_1605), .Z(n14_adj_821)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_229_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_457_i8_4_lut (.A(n6_adj_1408), .B(n14_adj_711), .C(n16331), 
         .D(n16345), .Z(n8_adj_496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_457_i8_4_lut.init = 16'hcfca;
    PFUMX PrioSelect_93_i16 (.BLUT(n11_adj_1497), .ALUT(n12_adj_1516), .C0(n16727), 
          .Z(n16_adj_1273)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_205_i14_3_lut_4_lut (.A(n22251), .B(n7762), .C(Z_N_387[0]), 
         .D(n10_adj_1604), .Z(n14_adj_973)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_205_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 PrioSelect_577_i13_3_lut_4_lut (.A(n22239), .B(n7908), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_1616)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_577_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_233_i14_3_lut_4_lut (.A(n22251), .B(n7762), .C(Z_N_387[7]), 
         .D(n10_adj_1603), .Z(n14_adj_639)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_233_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3146_3_lut_4_lut (.A(n22239), .B(n7908), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_1617)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i3146_3_lut_4_lut.init = 16'hf780;
    LUT4 i8911_2_lut_rep_681_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n10_adj_863), .D(n8_adj_708), .Z(n22248)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i8911_2_lut_rep_681_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_rep_571_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n11714), .D(n22279), .Z(n22138)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_571_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_595_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n7762), .D(n22279), .Z(n22162)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_595_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_619_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n16312), .D(n22279), .Z(n22186)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_619_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_691_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n10_adj_863), .D(n8_adj_708), .Z(n22258)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_691_3_lut_4_lut_4_lut.init = 16'h0008;
    PFUMX i18415 (.BLUT(n22323), .ALUT(n22324), .C0(instruction[15]), 
          .Z(n22325));
    PFUMX PrioSelect_89_i16 (.BLUT(n11_adj_1483), .ALUT(n12_adj_1515), .C0(n16727), 
          .Z(n16_adj_1272)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_541_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7908), .D(n22279), .Z(n22108)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_541_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 PrioSelect_245_i11_3_lut_4_lut (.A(n22255), .B(n7762), .C(instruction[2]), 
         .D(port_id_7__N_200[2]), .Z(n11_adj_1594)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_245_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_85_i16 (.BLUT(n11_adj_1472), .ALUT(n12_adj_1514), .C0(n16727), 
          .Z(n16_adj_1271)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_670_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n10_adj_863), .D(n8_adj_708), .Z(n22237)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_670_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_577_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n11714), .D(n22279), .Z(n22144)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_577_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_601_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n7762), .D(n22279), .Z(n22168)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_601_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX PrioSelect_81_i16 (.BLUT(n11_adj_1478), .ALUT(n12_adj_1517), .C0(n16727), 
          .Z(n16_adj_1270)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_625_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7876), 
         .C(n16312), .D(n22279), .Z(n22192)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_625_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i17618_2_lut_rep_558_3_lut_4_lut_4_lut_4_lut (.A(clk_in_c_enable_174), 
         .B(n22279), .C(n11778), .D(n11714), .Z(n22125)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i17618_2_lut_rep_558_3_lut_4_lut_4_lut_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_583_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7762), .D(n22279), .Z(n22150)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_583_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_643_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n7908), .D(n22279), .Z(n22210)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_643_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 PrioSelect_573_i13_3_lut_4_lut (.A(n22239), .B(n7908), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_1618)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_573_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_241_i11_3_lut_4_lut (.A(n22255), .B(n7762), .C(instruction[1]), 
         .D(port_id_7__N_200[1]), .Z(n11_adj_1597)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_241_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_249_i11_3_lut_4_lut (.A(n22255), .B(n7762), .C(instruction[3]), 
         .D(port_id_7__N_200[3]), .Z(n11_adj_1590)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_249_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_607_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n11778), 
         .C(n16312), .D(n22279), .Z(n22174)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_607_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i17580_4_lut (.A(n22141), .B(n22140), .C(n22138), .D(n17164), 
         .Z(n20182)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17580_4_lut.init = 16'hefee;
    LUT4 i13994_4_lut (.A(n22137), .B(n22136), .C(n213[2]), .D(n20955), 
         .Z(n17164)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i13994_4_lut.init = 16'h1011;
    L6MUX21 PrioSelect_585_i17 (.D0(n13_adj_1619), .D1(n16_adj_1620), .SD(n19570), 
            .Z(n17_adj_1399)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_565_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n11714), .D(n22279), .Z(n22132)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_565_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 PrioSelect_569_i13_3_lut_4_lut (.A(n22239), .B(n7908), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_1621)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_569_i13_3_lut_4_lut.init = 16'hf780;
    L6MUX21 PrioSelect_557_i17 (.D0(n13_adj_1622), .D1(n16_adj_1217), .SD(n19421), 
            .Z(n17_adj_1398)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17650_2_lut_3_lut_4_lut (.A(n22264), .B(n16392), .C(n20251), 
         .D(n7908), .Z(n19237)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17650_2_lut_3_lut_4_lut.init = 16'hf4f0;
    L6MUX21 PrioSelect_553_i17 (.D0(n13_adj_1623), .D1(n16_adj_1624), .SD(n19386), 
            .Z(n17_adj_1397)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_565_i13_3_lut_4_lut (.A(n22239), .B(n7908), .C(n703[2]), 
         .D(Z_N_378[2]), .Z(n13_adj_1625)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_565_i13_3_lut_4_lut.init = 16'hf780;
    L6MUX21 PrioSelect_525_i17 (.D0(n13_adj_1626), .D1(n16_adj_986), .SD(n19237), 
            .Z(n17_adj_1395)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 PrioSelect_521_i17 (.D0(n13_adj_1627), .D1(n16_adj_1628), .SD(n19202), 
            .Z(n17_adj_1393)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 PrioSelect_493_i17 (.D0(n13_adj_1629), .D1(n16_adj_988), .SD(n19053), 
            .Z(n17_adj_1391)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_253_i11_3_lut_4_lut (.A(n22255), .B(n7762), .C(instruction[4]), 
         .D(port_id_7__N_200[4]), .Z(n11_adj_1587)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_253_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_257_i11_3_lut_4_lut (.A(n22255), .B(n7762), .C(instruction[5]), 
         .D(port_id_7__N_200[5]), .Z(n11_adj_1480)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_257_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX i105 (.BLUT(n63_adj_1041), .ALUT(n14428), .C0(instruction[17]), 
          .Z(n105));
    LUT4 PrioSelect_261_i11_3_lut_4_lut (.A(n22255), .B(n7762), .C(instruction[6]), 
         .D(port_id_7__N_200[6]), .Z(n11_adj_1476)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(237[36:40])
    defparam PrioSelect_261_i11_3_lut_4_lut.init = 16'hf780;
    L6MUX21 PrioSelect_489_i17 (.D0(n13_adj_1630), .D1(n16), .SD(n19018), 
            .Z(n17_adj_1389)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_rep_589_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7762), .D(n22279), .Z(n22156)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_589_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 PrioSelect_265_i11_3_lut_4_lut (.A(n22253), .B(n7762), .C(Z_N_367[7]), 
         .D(instruction[7]), .Z(n11_adj_1631)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_265_i11_3_lut_4_lut.init = 16'hf780;
    L6MUX21 i16418 (.D0(n19584), .D1(n19585), .SD(instruction[6]), .Z(n19588));
    L6MUX21 i16419 (.D0(n19586), .D1(n19587), .SD(instruction[6]), .Z(n19589));
    L6MUX21 i16433 (.D0(n19599), .D1(n19600), .SD(instruction[6]), .Z(n19603));
    L6MUX21 PrioSelect_461_i17 (.D0(n13_adj_1632), .D1(n16_adj_953), .SD(n18869), 
            .Z(n17_adj_1388)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16434 (.D0(n19601), .D1(n19602), .SD(instruction[6]), .Z(n19604));
    L6MUX21 PrioSelect_457_i17 (.D0(n13_adj_497), .D1(n16_adj_493), .SD(n18834), 
            .Z(n17_adj_1386)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16448 (.D0(n19614), .D1(n19615), .SD(instruction[6]), .Z(n19618));
    L6MUX21 PrioSelect_429_i17 (.D0(n13_adj_1633), .D1(n16_adj_1026), .SD(n18685), 
            .Z(n17_adj_1385)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 PrioSelect_425_i17 (.D0(n13_adj_1634), .D1(n16_adj_514), .SD(n18650), 
            .Z(n17_adj_1382)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16449 (.D0(n19616), .D1(n19617), .SD(instruction[6]), .Z(n19619));
    L6MUX21 i16463 (.D0(n19629), .D1(n19630), .SD(instruction[6]), .Z(n19633));
    L6MUX21 i16464 (.D0(n19631), .D1(n19632), .SD(instruction[6]), .Z(n19634));
    L6MUX21 PrioSelect_397_i17 (.D0(n13_adj_1635), .D1(n16_adj_962), .SD(n18501), 
            .Z(n17_adj_1381)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16478 (.D0(n19644), .D1(n19645), .SD(instruction[6]), .Z(n19648));
    L6MUX21 PrioSelect_393_i17 (.D0(n13_adj_545), .D1(n16_adj_541), .SD(n18466), 
            .Z(n17_adj_1379)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16479 (.D0(n19646), .D1(n19647), .SD(instruction[6]), .Z(n19649));
    L6MUX21 i16493 (.D0(n19659), .D1(n19660), .SD(instruction[6]), .Z(n19663));
    LUT4 i17588_2_lut_3_lut_4_lut (.A(n22264), .B(n16392), .C(n20189), 
         .D(n7908), .Z(n19386)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17588_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 PrioSelect_237_i11_3_lut_4_lut (.A(n22253), .B(n7762), .C(Z_N_367[0]), 
         .D(instruction[0]), .Z(n11_adj_1636)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(263[50:54])
    defparam PrioSelect_237_i11_3_lut_4_lut.init = 16'hf780;
    L6MUX21 i16494 (.D0(n19661), .D1(n19662), .SD(instruction[6]), .Z(n19664));
    L6MUX21 PrioSelect_365_i17 (.D0(n13_adj_1637), .D1(n16_adj_1084), .SD(n18317), 
            .Z(n17_adj_1378)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16508 (.D0(n19674), .D1(n19675), .SD(instruction[6]), .Z(n19678));
    L6MUX21 i16509 (.D0(n19676), .D1(n19677), .SD(instruction[6]), .Z(n19679));
    L6MUX21 PrioSelect_361_i17 (.D0(n13_adj_1638), .D1(n16_adj_560), .SD(n18282), 
            .Z(n17_adj_1376)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16612 (.D0(n19778), .D1(n19779), .SD(instruction[6]), .Z(n19782));
    L6MUX21 PrioSelect_333_i17 (.D0(n13_adj_1639), .D1(n16_adj_967), .SD(n18133), 
            .Z(n17_adj_1374)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16613 (.D0(n19780), .D1(n19781), .SD(instruction[6]), .Z(n19783));
    PFUMX i16414 (.BLUT(n19576), .ALUT(n19577), .C0(instruction[5]), .Z(n19584));
    PFUMX i16415 (.BLUT(n19578), .ALUT(n19579), .C0(instruction[5]), .Z(n19585));
    L6MUX21 PrioSelect_329_i17 (.D0(n13_adj_579), .D1(n16_adj_576), .SD(n18098), 
            .Z(n17_adj_1373)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 PrioSelect_301_i17 (.D0(n13_adj_1640), .D1(n16_adj_1132), .SD(n17949), 
            .Z(n17_adj_1372)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 PrioSelect_297_i17 (.D0(n13_adj_1641), .D1(n16_adj_599), .SD(n17914), 
            .Z(n17_adj_1370)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 PrioSelect_269_i17 (.D0(n13_adj_1642), .D1(n16_adj_969), .SD(n17765), 
            .Z(n17_adj_1369)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16416 (.BLUT(n19580), .ALUT(n19581), .C0(instruction[5]), .Z(n19586));
    L6MUX21 PrioSelect_265_i17 (.D0(n13_adj_619), .D1(n16_adj_616), .SD(n17730), 
            .Z(n17_adj_1368)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16417 (.BLUT(n19582), .ALUT(n19583), .C0(instruction[5]), .Z(n19587));
    LUT4 i17596_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n16392), .C(n11714), 
         .D(n22263), .Z(n17155)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17596_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h040c;
    PFUMX i16429 (.BLUT(n19591), .ALUT(n19592), .C0(instruction[5]), .Z(n19599));
    L6MUX21 PrioSelect_237_i17 (.D0(n13_adj_1643), .D1(n16_adj_1143), .SD(n17581), 
            .Z(n17_adj_1367)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 PrioSelect_233_i17 (.D0(n13_adj_1644), .D1(n16_adj_641), .SD(n17546), 
            .Z(n17_adj_1366)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17698_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n22258), .B(n7762), .C(n22255), 
         .D(n22253), .Z(n17722)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam i17698_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hccc8;
    L6MUX21 PrioSelect_205_i17 (.D0(n13_adj_1645), .D1(n16_adj_975), .SD(n17397), 
            .Z(n17_adj_1361)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16430 (.BLUT(n19593), .ALUT(n19594), .C0(instruction[5]), .Z(n19600));
    LUT4 PrioSelect_237_i12_3_lut_4_lut (.A(n22258), .B(n7762), .C(Z_N_378[0]), 
         .D(n11_adj_1636), .Z(n12_adj_1646)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_237_i12_3_lut_4_lut.init = 16'hf780;
    PFUMX i16431 (.BLUT(n19595), .ALUT(n19596), .C0(instruction[5]), .Z(n19601));
    L6MUX21 PrioSelect_201_i17 (.D0(n13_adj_675), .D1(n16_adj_671), .SD(n17362), 
            .Z(n17_adj_1360)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_265_i12_3_lut_4_lut (.A(n22258), .B(n7762), .C(Z_N_378[7]), 
         .D(n11_adj_1631), .Z(n12_adj_618)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(275[49:53])
    defparam PrioSelect_265_i12_3_lut_4_lut.init = 16'hf780;
    L6MUX21 PrioSelect_173_i17 (.D0(n13_adj_1647), .D1(n16_adj_1163), .SD(n17213), 
            .Z(n17_adj_1648)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_561_i13_3_lut_4_lut (.A(n22239), .B(n7908), .C(n703[1]), 
         .D(Z_N_378[1]), .Z(n13_adj_1649)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_561_i13_3_lut_4_lut.init = 16'hf780;
    L6MUX21 PrioSelect_169_i17 (.D0(n13_adj_1650), .D1(n16_adj_756), .SD(n17178), 
            .Z(n17_adj_1651)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16432 (.BLUT(n19597), .ALUT(n19598), .C0(instruction[5]), .Z(n19602));
    L6MUX21 PrioSelect_141_i17 (.D0(n13_adj_1652), .D1(n16_adj_980), .SD(n17029), 
            .Z(n17_adj_1613)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 PrioSelect_137_i17 (.D0(n13_adj_847), .D1(n16_adj_842), .SD(n16994), 
            .Z(n17_adj_1611)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16444 (.BLUT(n19606), .ALUT(n19607), .C0(instruction[5]), .Z(n19614));
    L6MUX21 PrioSelect_109_i17 (.D0(n13_adj_1653), .D1(n16_adj_1182), .SD(n16845), 
            .Z(n17_adj_1593)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 PrioSelect_105_i17 (.D0(n13_adj_1654), .D1(n16_adj_879), .SD(n16810), 
            .Z(n17_adj_1592)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16445 (.BLUT(n19608), .ALUT(n19609), .C0(instruction[5]), .Z(n19615));
    L6MUX21 PrioSelect_77_i17 (.D0(n13_adj_1655), .D1(n16_adj_983), .SD(n16662), 
            .Z(n17_adj_1513)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16446 (.BLUT(n19610), .ALUT(n19611), .C0(instruction[5]), .Z(n19616));
    PFUMX i16447 (.BLUT(n19612), .ALUT(n19613), .C0(instruction[5]), .Z(n19617));
    L6MUX21 i116 (.D0(n58), .D1(n85), .SD(n16618), .Z(n64_adj_1492));
    LUT4 PrioSelect_241_i12_3_lut_4_lut (.A(n22254), .B(n7762), .C(n1108[1]), 
         .D(Z_N_367[1]), .Z(n12_adj_1598)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_241_i12_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_557_i13 (.BLUT(n4_adj_1020), .ALUT(n12_adj_1578), .C0(n19562), 
          .Z(n13_adj_1622)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16459 (.BLUT(n19621), .ALUT(n19622), .C0(instruction[5]), .Z(n19629));
    PFUMX i16460 (.BLUT(n19623), .ALUT(n19624), .C0(instruction[5]), .Z(n19630));
    LUT4 i17581_2_lut_3_lut_4_lut (.A(n22264), .B(n16392), .C(n20182), 
         .D(n11714), .Z(n17178)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17581_2_lut_3_lut_4_lut.init = 16'hf0f4;
    PFUMX PrioSelect_525_i13 (.BLUT(n4_adj_1016), .ALUT(n12_adj_1570), .C0(n19378), 
          .Z(n13_adj_1626)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16461 (.BLUT(n19625), .ALUT(n19626), .C0(instruction[5]), .Z(n19631));
    LUT4 PrioSelect_245_i12_3_lut_4_lut (.A(n22254), .B(n7762), .C(n1108[2]), 
         .D(Z_N_367[2]), .Z(n12_adj_1595)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_245_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_613_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n16312), .D(n22279), .Z(n22180)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_613_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX i16462 (.BLUT(n19627), .ALUT(n19628), .C0(instruction[5]), .Z(n19632));
    PFUMX PrioSelect_493_i13 (.BLUT(n4_adj_1012), .ALUT(n12_adj_1518), .C0(n19194), 
          .Z(n13_adj_1629)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i1_2_lut_adj_202 (.A(instruction[9]), .B(instruction[8]), .Z(n16392)) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(219[39:43])
    defparam i1_2_lut_adj_202.init = 16'h2222;
    LUT4 PrioSelect_249_i12_3_lut_4_lut (.A(n22254), .B(n7762), .C(n1108[3]), 
         .D(Z_N_367[3]), .Z(n12_adj_1591)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_249_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_253_i12_3_lut_4_lut (.A(n22254), .B(n7762), .C(n1108[4]), 
         .D(Z_N_367[4]), .Z(n12_adj_1588)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_253_i12_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_489_i13 (.BLUT(n8_adj_996), .ALUT(n12_adj_1427), .C0(n19010), 
          .Z(n13_adj_1630)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16474 (.BLUT(n19636), .ALUT(n19637), .C0(instruction[5]), .Z(n19644));
    LUT4 i1_2_lut_rep_650_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n7726), 
         .C(n7908), .D(n22279), .Z(n22217)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_650_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_664_3_lut_4_lut_4_lut (.A(clk_in_c_enable_174), .B(n16392), 
         .C(n10_adj_863), .D(n8_adj_708), .Z(n22231)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_664_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 PrioSelect_585_i10_3_lut_4_lut (.A(n22239), .B(n7908), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_1656)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_585_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i17672_4_lut_4_lut (.A(clk_in_c_enable_109), .B(n8050), .C(n10_adj_812), 
         .D(n22300), .Z(clk_in_c_enable_113)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i17672_4_lut_4_lut.init = 16'h0002;
    LUT4 i17688_2_lut_3_lut_4_lut (.A(n22264), .B(n16392), .C(n20289), 
         .D(n11714), .Z(n17029)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17688_2_lut_3_lut_4_lut.init = 16'hf0f4;
    LUT4 i17687_4_lut (.A(n22141), .B(n22140), .C(n22138), .D(n17011), 
         .Z(n20289)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17687_4_lut.init = 16'hefee;
    PFUMX PrioSelect_461_i13 (.BLUT(n4_adj_992), .ALUT(n12_adj_1428), .C0(n19010), 
          .Z(n13_adj_1632)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_257_i12_3_lut_4_lut (.A(n22254), .B(n7762), .C(n1108[5]), 
         .D(Z_N_367[5]), .Z(n12_adj_1481)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_257_i12_3_lut_4_lut.init = 16'hf780;
    PFUMX i16475 (.BLUT(n19638), .ALUT(n19639), .C0(instruction[5]), .Z(n19645));
    LUT4 PrioSelect_169_i19_4_lut (.A(n17_adj_1651), .B(in_port[7]), .C(n22104), 
         .D(n346[2]), .Z(n491)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_169_i19_4_lut.init = 16'hc0ca;
    LUT4 i17655_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n16392), .C(n7762), 
         .D(n22263), .Z(n17891)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17655_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i17630_2_lut_3_lut_4_lut (.A(n22264), .B(n16392), .C(n20231), 
         .D(n7762), .Z(n17914)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17630_2_lut_3_lut_4_lut.init = 16'hf4f0;
    PFUMX i16476 (.BLUT(n19640), .ALUT(n19641), .C0(instruction[5]), .Z(n19646));
    PFUMX i18413 (.BLUT(n22320), .ALUT(n22321), .C0(instruction[16]), 
          .Z(n22322));
    LUT4 i17763_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n16392), .C(n16312), 
         .D(n22263), .Z(n18627)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17763_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    LUT4 i17686_2_lut_3_lut_4_lut (.A(n22264), .B(n16392), .C(n20287), 
         .D(n7762), .Z(n17765)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17686_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 PrioSelect_561_i14_3_lut_4_lut (.A(n22240), .B(n7908), .C(Z_N_387[1]), 
         .D(n13_adj_1649), .Z(n14_adj_1093)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_561_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i13841_4_lut (.A(n22137), .B(n22136), .C(n213[2]), .D(n17002), 
         .Z(n17011)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i13841_4_lut.init = 16'h1011;
    LUT4 PrioSelect_261_i12_3_lut_4_lut (.A(n22254), .B(n7762), .C(n1108[6]), 
         .D(Z_N_367[6]), .Z(n12_adj_1477)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_261_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_237_i15_3_lut_4_lut (.A(n22254), .B(n7762), .C(n1108[0]), 
         .D(n5_adj_1183), .Z(n15_adj_1142)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_237_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_565_i14_3_lut_4_lut (.A(n22240), .B(n7908), .C(Z_N_387[2]), 
         .D(n13_adj_1625), .Z(n14_adj_1110)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_565_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17760_2_lut_3_lut_4_lut (.A(n22264), .B(n16392), .C(n20361), 
         .D(n16312), .Z(n18650)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17760_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i17776_2_lut_3_lut_4_lut (.A(n22264), .B(n16392), .C(n20377), 
         .D(n16312), .Z(n18501)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17776_2_lut_3_lut_4_lut.init = 16'hf4f0;
    PFUMX PrioSelect_429_i13 (.BLUT(n4_adj_972), .ALUT(n12_adj_1267), .C0(n18826), 
          .Z(n13_adj_1633)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_265_i15_3_lut_4_lut (.A(n22254), .B(n7762), .C(n1108[7]), 
         .D(n9_adj_876), .Z(n15_adj_615)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam PrioSelect_265_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_569_i14_3_lut_4_lut (.A(n22240), .B(n7908), .C(Z_N_387[3]), 
         .D(n13_adj_1621), .Z(n14_adj_1101)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_569_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 PrioSelect_265_i10_3_lut_4_lut (.A(n22259), .B(n7762), .C(n703[7]), 
         .D(port_id_7__N_200[7]), .Z(n10_adj_735)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_265_i10_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_425_i13 (.BLUT(n8_adj_959), .ALUT(n12_adj_1231), .C0(n18642), 
          .Z(n13_adj_1634)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 i17591_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n22264), .B(n16392), .C(n7908), 
         .D(n22263), .Z(n19363)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(369[51:55])
    defparam i17591_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h40c0;
    PFUMX PrioSelect_397_i13 (.BLUT(n4_adj_950), .ALUT(n12_adj_1232), .C0(n18642), 
          .Z(n13_adj_1635)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_573_i14_3_lut_4_lut (.A(n22240), .B(n7908), .C(Z_N_387[4]), 
         .D(n13_adj_1618), .Z(n14_adj_1098)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_573_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX i16477 (.BLUT(n19642), .ALUT(n19643), .C0(instruction[5]), .Z(n19647));
    PFUMX i16489 (.BLUT(n19651), .ALUT(n19652), .C0(instruction[5]), .Z(n19659));
    PFUMX i16490 (.BLUT(n19653), .ALUT(n19654), .C0(instruction[5]), .Z(n19660));
    PFUMX i16491 (.BLUT(n19655), .ALUT(n19656), .C0(instruction[5]), .Z(n19661));
    LUT4 PrioSelect_173_i19_4_lut (.A(n17_adj_1648), .B(in_port[0]), .C(n22103), 
         .D(n346[3]), .Z(n495)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam PrioSelect_173_i19_4_lut.init = 16'hc0ca;
    PFUMX PrioSelect_365_i13 (.BLUT(n4_adj_948), .ALUT(n12_adj_1196), .C0(n18306), 
          .Z(n13_adj_1637)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16492 (.BLUT(n19657), .ALUT(n19658), .C0(instruction[5]), .Z(n19662));
    PFUMX i16504 (.BLUT(n19666), .ALUT(n19667), .C0(instruction[5]), .Z(n19674));
    PFUMX i16505 (.BLUT(n19668), .ALUT(n19669), .C0(instruction[5]), .Z(n19675));
    LUT4 i1059_3_lut_4_lut (.A(st[2]), .B(n22305), .C(st[3]), .D(st[4]), 
         .Z(stack_N_397[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(203[23:27])
    defparam i1059_3_lut_4_lut.init = 16'h7f80;
    PFUMX PrioSelect_361_i13 (.BLUT(n8_adj_946), .ALUT(n12_adj_1146), .C0(n18274), 
          .Z(n13_adj_1638)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16506 (.BLUT(n19670), .ALUT(n19671), .C0(instruction[5]), .Z(n19676));
    LUT4 PrioSelect_557_i14_3_lut_4_lut (.A(n22240), .B(n7908), .C(Z_N_387[0]), 
         .D(n10_adj_1617), .Z(n14_adj_1215)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_557_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX i16507 (.BLUT(n19672), .ALUT(n19673), .C0(instruction[5]), .Z(n19677));
    PFUMX i16515 (.BLUT(n19681), .ALUT(n19682), .C0(instruction[9]), .Z(n19685));
    PFUMX PrioSelect_333_i13 (.BLUT(n4_adj_942), .ALUT(n12_adj_1147), .C0(n18274), 
          .Z(n13_adj_1639)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16516 (.BLUT(n19683), .ALUT(n19684), .C0(instruction[9]), .Z(n19686));
    LUT4 PrioSelect_577_i14_3_lut_4_lut (.A(n22240), .B(n7908), .C(Z_N_387[5]), 
         .D(n13_adj_1616), .Z(n14_adj_1105)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_577_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_301_i13 (.BLUT(n4_adj_939), .ALUT(n12_adj_1052), .C0(n18090), 
          .Z(n13_adj_1640)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16522 (.BLUT(n19688), .ALUT(n19689), .C0(instruction[9]), .Z(n19692));
    PFUMX i16523 (.BLUT(n19690), .ALUT(n19691), .C0(instruction[9]), .Z(n19693));
    LUT4 PrioSelect_581_i14_3_lut_4_lut (.A(n22240), .B(n7908), .C(Z_N_387[6]), 
         .D(n13_adj_1615), .Z(n14_adj_1088)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_581_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_297_i13 (.BLUT(n8_adj_936), .ALUT(n12_adj_859), .C0(n17906), 
          .Z(n13_adj_1641)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16529 (.BLUT(n19695), .ALUT(n19696), .C0(instruction[9]), .Z(n19699));
    PFUMX i16530 (.BLUT(n19697), .ALUT(n19698), .C0(instruction[9]), .Z(n19700));
    LUT4 i8711_2_lut_rep_718_3_lut_3_lut_4_lut (.A(st_zc[2]), .B(n22306), 
         .C(st_zc[3]), .D(st_zc[4]), .Z(n22285)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(206[26:38])
    defparam i8711_2_lut_rep_718_3_lut_3_lut_4_lut.init = 16'h7ff8;
    LUT4 i17700_4_lut (.A(n22135), .B(n22134), .C(n22132), .D(n16980), 
         .Z(n20302)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17700_4_lut.init = 16'hefee;
    LUT4 i1_2_lut_rep_715_3_lut_3_lut_4_lut (.A(st_zc[2]), .B(n22306), .C(st_zc[3]), 
         .D(st_zc[4]), .Z(n22282)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(206[26:38])
    defparam i1_2_lut_rep_715_3_lut_3_lut_4_lut.init = 16'h0078;
    LUT4 i13810_4_lut (.A(n22131), .B(n22130), .C(n213[1]), .D(n20914), 
         .Z(n16980)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i13810_4_lut.init = 16'h1011;
    LUT4 i1095_3_lut_rep_720_4_lut (.A(st_zc[2]), .B(n22306), .C(st_zc[3]), 
         .D(st_zc[4]), .Z(n22287)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(206[26:38])
    defparam i1095_3_lut_rep_720_4_lut.init = 16'h7f80;
    PFUMX PrioSelect_269_i13 (.BLUT(n4_adj_928), .ALUT(n12_adj_860), .C0(n17906), 
          .Z(n13_adj_1642)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_585_i14_3_lut_4_lut (.A(n22240), .B(n7908), .C(Z_N_387[7]), 
         .D(n10_adj_1656), .Z(n14_adj_1657)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(333[49:53])
    defparam PrioSelect_585_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX i16536 (.BLUT(n19702), .ALUT(n19703), .C0(instruction[9]), .Z(n19706));
    LUT4 i2026_3_lut_4_lut (.A(n22259), .B(n7762), .C(n703[0]), .D(port_id_7__N_200[0]), 
         .Z(n10_adj_733)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i2026_3_lut_4_lut.init = 16'hf780;
    PFUMX i16537 (.BLUT(n19704), .ALUT(n19705), .C0(instruction[9]), .Z(n19707));
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(st_zc[2]), .B(n22306), .C(st_zc[3]), 
         .D(st_zc[4]), .Z(n7746)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(206[26:38])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h0780;
    PFUMX PrioSelect_237_i13 (.BLUT(n4_adj_923), .ALUT(n12_adj_1646), .C0(n17722), 
          .Z(n13_adj_1643)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_261_i13_3_lut_4_lut (.A(n22259), .B(n7762), .C(n703[6]), 
         .D(Z_N_378[6]), .Z(n13_adj_725)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_261_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i17741_3_lut_rep_729 (.A(jp), .B(rst_n_in), .C(clk_in_c_enable_109), 
         .Z(clk_in_c_enable_174)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i17741_3_lut_rep_729.init = 16'h4040;
    LUT4 i1_2_lut_rep_713_4_lut (.A(jp), .B(rst_n_in), .C(clk_in_c_enable_109), 
         .D(n16392), .Z(n22280)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_rep_713_4_lut.init = 16'h4000;
    LUT4 i17773_4_lut (.A(n22135), .B(n22134), .C(n22132), .D(n16827), 
         .Z(n20375)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i17773_4_lut.init = 16'hefee;
    LUT4 PrioSelect_257_i13_3_lut_4_lut (.A(n22259), .B(n7762), .C(n703[5]), 
         .D(Z_N_378[5]), .Z(n13_adj_717)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_257_i13_3_lut_4_lut.init = 16'hf780;
    PFUMX i16543 (.BLUT(n19709), .ALUT(n19710), .C0(instruction[9]), .Z(n19713));
    PFUMX PrioSelect_233_i13 (.BLUT(n8_adj_915), .ALUT(n12_adj_1586), .C0(n17538), 
          .Z(n13_adj_1644)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16544 (.BLUT(n19711), .ALUT(n19712), .C0(instruction[9]), .Z(n19714));
    LUT4 i1_2_lut_adj_203 (.A(instruction[8]), .B(instruction[9]), .Z(n7876)) /* synthesis lut_function=(A (B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(228[39:43])
    defparam i1_2_lut_adj_203.init = 16'h8888;
    PFUMX PrioSelect_205_i13 (.BLUT(n4_adj_902), .ALUT(n12_adj_1589), .C0(n17538), 
          .Z(n13_adj_1645)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_253_i13_3_lut_4_lut (.A(n22259), .B(n7762), .C(n703[4]), 
         .D(Z_N_378[4]), .Z(n13_adj_714)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_253_i13_3_lut_4_lut.init = 16'hf780;
    PFUMX i16550 (.BLUT(n19716), .ALUT(n19717), .C0(instruction[9]), .Z(n19720));
    PFUMX PrioSelect_173_i13 (.BLUT(n4_adj_892), .ALUT(n12_adj_814), .C0(n17354), 
          .Z(n13_adj_1647)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16551 (.BLUT(n19718), .ALUT(n19719), .C0(instruction[9]), .Z(n19721));
    LUT4 i13657_4_lut (.A(n22131), .B(n22130), .C(n213[1]), .D(n16818), 
         .Z(n16827)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(100[41:42])
    defparam i13657_4_lut.init = 16'h1011;
    PFUMX i16557 (.BLUT(n19723), .ALUT(n19724), .C0(instruction[9]), .Z(n19727));
    LUT4 PrioSelect_557_i5_3_lut_4_lut (.A(n22227), .B(n22281), .C(n13_adj_731), 
         .D(n14_adj_711), .Z(n5_adj_1612)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam PrioSelect_557_i5_3_lut_4_lut.init = 16'hf780;
    PFUMX i16558 (.BLUT(n19725), .ALUT(n19726), .C0(instruction[9]), .Z(n19728));
    LUT4 i13385_2_lut_rep_709_2_lut_4_lut (.A(jp), .B(rst_n_in), .C(clk_in_c_enable_109), 
         .D(n10_adj_698), .Z(n22276)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i13385_2_lut_rep_709_2_lut_4_lut.init = 16'hffbf;
    PFUMX i16564 (.BLUT(n19730), .ALUT(n19731), .C0(instruction[9]), .Z(n19734));
    PFUMX PrioSelect_169_i13 (.BLUT(n8_adj_885), .ALUT(n12_adj_1444), .C0(n17170), 
          .Z(n13_adj_1650)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16565 (.BLUT(n19732), .ALUT(n19733), .C0(instruction[9]), .Z(n19735));
    LUT4 i3242_3_lut_4_lut (.A(n22227), .B(n22281), .C(n13_adj_748), .D(n13_adj_744), 
         .Z(n10_adj_1089)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/top.v(59[13:24])
    defparam i3242_3_lut_4_lut.init = 16'hf780;
    PFUMX i16569 (.BLUT(n19737), .ALUT(n19738), .C0(instruction[9]), .Z(n13_adj_736));
    PFUMX PrioSelect_141_i13 (.BLUT(n4_adj_881), .ALUT(n12_adj_1447), .C0(n17170), 
          .Z(n13_adj_1652)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16572 (.BLUT(n19740), .ALUT(n19741), .C0(instruction[9]), .Z(n19742));
    PFUMX i16575 (.BLUT(n19743), .ALUT(n19744), .C0(instruction[9]), .Z(n13_adj_731));
    LUT4 i17599_2_lut_rep_518_3_lut_3_lut_4_lut_4_lut (.A(n22267), .B(n16392), 
         .C(n11714), .D(n22268), .Z(n22085)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((C)+!B))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam i17599_2_lut_rep_518_3_lut_3_lut_4_lut_4_lut.init = 16'h040c;
    LUT4 i1_2_lut_rep_710_2_lut_4_lut (.A(jp), .B(rst_n_in), .C(clk_in_c_enable_109), 
         .D(n8_adj_695), .Z(n22277)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_2_lut_rep_710_2_lut_4_lut.init = 16'hffbf;
    LUT4 i1448_2_lut_rep_731 (.A(st_zc[0]), .B(st_zc[1]), .Z(n22298)) /* synthesis lut_function=(A+(B)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(376[91:109])
    defparam i1448_2_lut_rep_731.init = 16'heeee;
    PFUMX i18411 (.BLUT(n22317), .ALUT(n22318), .C0(instruction[15]), 
          .Z(n22319));
    PFUMX PrioSelect_109_i13 (.BLUT(n4_adj_856), .ALUT(n12_adj_1317), .C0(n16986), 
          .Z(n13_adj_1653)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16578 (.BLUT(n19746), .ALUT(n19747), .C0(instruction[9]), .Z(n19748));
    LUT4 i1207_2_lut_3_lut_4_lut (.A(st_zc[0]), .B(st_zc[1]), .C(st_zc[3]), 
         .D(st_zc[2]), .Z(n8_adj_1453)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(376[91:109])
    defparam i1207_2_lut_3_lut_4_lut.init = 16'hfffe;
    PFUMX i16581 (.BLUT(n19749), .ALUT(n19750), .C0(instruction[9]), .Z(n13_adj_748));
    PFUMX i16584 (.BLUT(n19752), .ALUT(n19753), .C0(instruction[9]), .Z(n19754));
    PFUMX PrioSelect_105_i13 (.BLUT(n8_adj_853), .ALUT(n12_adj_1508), .C0(n16802), 
          .Z(n13_adj_1654)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16587 (.BLUT(n19755), .ALUT(n19756), .C0(instruction[9]), .Z(n13_adj_515));
    PFUMX i16590 (.BLUT(n19758), .ALUT(n19759), .C0(instruction[9]), .Z(n19760));
    PFUMX i16593 (.BLUT(n19761), .ALUT(n19762), .C0(instruction[9]), .Z(n13_adj_744));
    PFUMX i16596 (.BLUT(n19764), .ALUT(n19765), .C0(instruction[9]), .Z(n19766));
    PFUMX PrioSelect_77_i13 (.BLUT(n4_adj_850), .ALUT(n12_adj_1509), .C0(n16802), 
          .Z(n13_adj_1655)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16599 (.BLUT(n19767), .ALUT(n19768), .C0(instruction[9]), .Z(n13_adj_516));
    PFUMX i120 (.BLUT(n14780), .ALUT(n19), .C0(instruction[14]), .Z(n58));
    PFUMX i16608 (.BLUT(n19770), .ALUT(n19771), .C0(instruction[5]), .Z(n19778));
    PFUMX i16609 (.BLUT(n19772), .ALUT(n19773), .C0(instruction[5]), .Z(n19779));
    PFUMX i16610 (.BLUT(n19774), .ALUT(n19775), .C0(instruction[5]), .Z(n19780));
    PFUMX i16611 (.BLUT(n19776), .ALUT(n19777), .C0(instruction[5]), .Z(n19781));
    PFUMX i16617 (.BLUT(n19785), .ALUT(n19786), .C0(instruction[9]), .Z(n19787));
    PFUMX i109 (.BLUT(n14803), .ALUT(n16391), .C0(instruction[13]), .Z(n53));
    PFUMX i16620 (.BLUT(n19788), .ALUT(n19789), .C0(instruction[9]), .Z(n13_adj_739));
    PFUMX i16623 (.BLUT(n19791), .ALUT(n19792), .C0(instruction[9]), .Z(n19793));
    PFUMX i16626 (.BLUT(n19794), .ALUT(n19795), .C0(instruction[9]), .Z(n19796));
    PFUMX i16629 (.BLUT(n19797), .ALUT(n19798), .C0(instruction[9]), .Z(n5_adj_737));
    PFUMX PrioSelect_585_i16 (.BLUT(n14_adj_1657), .ALUT(n15_adj_1614), 
          .C0(n19574), .Z(n16_adj_1620)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16776 (.D0(n19944), .D1(n19945), .SD(st_zc[3]), .Z(n19946));
    L6MUX21 i16791 (.D0(n19959), .D1(n19960), .SD(st_zc[3]), .Z(n19961));
    PFUMX PrioSelect_585_i13 (.BLUT(n8_adj_839), .ALUT(n12_adj_1580), .C0(n19562), 
          .Z(n13_adj_1619)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16774 (.D0(n19940), .D1(n19941), .SD(st_zc[2]), .Z(n19944));
    L6MUX21 i16775 (.D0(n19942), .D1(n19943), .SD(st_zc[2]), .Z(n19945));
    L6MUX21 i16789 (.D0(n19955), .D1(n19956), .SD(st_zc[2]), .Z(n19959));
    L6MUX21 i16790 (.D0(n19957), .D1(n19958), .SD(st_zc[2]), .Z(n19960));
    PFUMX PrioSelect_581_i19 (.BLUT(n15_adj_1090), .ALUT(n17_adj_1120), 
          .C0(n19545), .Z(n922)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_577_i19 (.BLUT(n15_adj_1106), .ALUT(n17_adj_1118), 
          .C0(n19545), .Z(n918)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_573_i19 (.BLUT(n15_adj_1099), .ALUT(n17_adj_1115), 
          .C0(n19545), .Z(n914)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_569_i19 (.BLUT(n15_adj_1102), .ALUT(n17_adj_1113), 
          .C0(n19545), .Z(n910)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_565_i19 (.BLUT(n15_adj_1111), .ALUT(n17_adj_1109), 
          .C0(n19545), .Z(n906)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_561_i19 (.BLUT(n15_adj_1095), .ALUT(n17_adj_1104), 
          .C0(n19545), .Z(n902)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_553_i16 (.BLUT(n14_adj_1199), .ALUT(n15_adj_1176), 
          .C0(n19390), .Z(n16_adj_1624)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_553_i13 (.BLUT(n8_adj_782), .ALUT(n12_adj_1572), .C0(n19378), 
          .Z(n13_adj_1623)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i18409 (.BLUT(n22314), .ALUT(n22315), .C0(st_zc[3]), .Z(n22316));
    LUT4 i8590_2_lut_3_lut (.A(st_zc[0]), .B(st_zc[1]), .C(stack_zc_20_1), 
         .Z(n21)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(376[91:109])
    defparam i8590_2_lut_3_lut.init = 16'h1010;
    PFUMX PrioSelect_549_i19 (.BLUT(n15_adj_1060), .ALUT(n17_adj_1310), 
          .C0(n19361), .Z(n890)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    LUT4 PrioSelect_249_i13_3_lut_4_lut (.A(n22259), .B(n7762), .C(n703[3]), 
         .D(Z_N_378[3]), .Z(n13_adj_703)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // f:/home/mini-mcu/step_fpga/mcu.v(281[53:57])
    defparam PrioSelect_249_i13_3_lut_4_lut.init = 16'hf780;
    PFUMX PrioSelect_545_i19 (.BLUT(n15_adj_1081), .ALUT(n17_adj_1308), 
          .C0(n19361), .Z(n886)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_541_i19 (.BLUT(n15_adj_1069), .ALUT(n17_adj_1306), 
          .C0(n19361), .Z(n882)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_537_i19 (.BLUT(n15_adj_1078), .ALUT(n17_adj_1302), 
          .C0(n19361), .Z(n878)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_533_i19 (.BLUT(n15_adj_1087), .ALUT(n17_adj_1300), 
          .C0(n19361), .Z(n874)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX PrioSelect_529_i19 (.BLUT(n15_adj_1063), .ALUT(n17_adj_1298), 
          .C0(n19361), .Z(n870)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16517 (.D0(n19685), .D1(n19686), .SD(instruction[10]), .Z(n7_adj_481));
    PFUMX PrioSelect_521_i16 (.BLUT(n14_adj_1549), .ALUT(n15_adj_632), .C0(n19206), 
          .Z(n16_adj_1628)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    L6MUX21 i16524 (.D0(n19692), .D1(n19693), .SD(instruction[10]), .Z(n7_adj_479));
    PFUMX PrioSelect_521_i13 (.BLUT(n8_adj_722), .ALUT(n12_adj_1519), .C0(n19194), 
          .Z(n13_adj_1627)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16758 (.BLUT(n19926), .ALUT(n19927), .C0(st_zc[1]), .Z(n19928));
    PFUMX i16761 (.BLUT(n19929), .ALUT(n19930), .C0(st_zc[1]), .Z(n19931));
    PFUMX PrioSelect_517_i19 (.BLUT(n15_adj_1505), .ALUT(n17_adj_1242), 
          .C0(n19177), .Z(n858)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16770 (.BLUT(n19932), .ALUT(n19933), .C0(st_zc[1]), .Z(n19940));
    PFUMX PrioSelect_513_i19 (.BLUT(n15_adj_1511), .ALUT(n17_adj_1238), 
          .C0(n19177), .Z(n854)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16771 (.BLUT(n19934), .ALUT(n19935), .C0(st_zc[1]), .Z(n19941));
    PFUMX i16772 (.BLUT(n19936), .ALUT(n19937), .C0(st_zc[1]), .Z(n19942));
    PFUMX PrioSelect_509_i19 (.BLUT(n15_adj_1521), .ALUT(n17_adj_1236), 
          .C0(n19177), .Z(n850)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16773 (.BLUT(n19938), .ALUT(n19939), .C0(st_zc[1]), .Z(n19943));
    PFUMX i16785 (.BLUT(n19947), .ALUT(n19948), .C0(st_zc[1]), .Z(n19955));
    PFUMX i16786 (.BLUT(n19949), .ALUT(n19950), .C0(st_zc[1]), .Z(n19956));
    PFUMX PrioSelect_505_i19 (.BLUT(n15_adj_495), .ALUT(n17_adj_1234), .C0(n19177), 
          .Z(n846)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    PFUMX i16787 (.BLUT(n19951), .ALUT(n19952), .C0(st_zc[1]), .Z(n19957));
    PFUMX i16788 (.BLUT(n19953), .ALUT(n19954), .C0(st_zc[1]), .Z(n19958));
    PFUMX PrioSelect_501_i19 (.BLUT(n15_adj_530), .ALUT(n17_adj_1230), .C0(n19177), 
          .Z(n842)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=2, LSE_LLINE=90, LSE_RLINE=102 */ ;
    
endmodule
