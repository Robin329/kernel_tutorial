always @(posedge clk or negedge rst)
begin
   if(rst==1'b0)begin

   end
   else begin

   end 
end