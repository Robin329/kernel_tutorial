`timescale 1ns / 1ps

module rom(
    input          clk,
    input [11:0]address,       //程序取址地址
    output[17:0]instruction,   //指令输入
    input       enable   //程序rom使能 1-->使能
);
(* ram_style="distributed" *)reg [17:0] y/* synthesis syn_ramstyle = "block_ram" */;
assign instruction = y;
always@(posedge clk) begin
    if(enable)begin
      case(address)
            12'd0 : y <= 18'h01AFE ;
            12'd1 : y <= 18'h2DA01 ;
            12'd2 : y <= 18'h2FA01 ;
            12'd3 : y <= 18'h01B66 ;
            12'd4 : y <= 18'h2FB00 ;
            12'd5 : y <= 18'h2DB00 ;
            12'd6 : y <= 18'h01C07 ;
            12'd7 : y <= 18'h2DC02 ;
            12'd8 : y <= 18'h09D00 ;
            12'd9 : y <= 18'h28001 ;
            12'd10 : y <= 18'h09D00 ;
            12'd11 : y <= 18'h14D06 ;
            12'd12 : y <= 18'h3E029 ;
            12'd13 : y <= 18'h14D06 ;
            12'd14 : y <= 18'h3E022 ;
            12'd15 : y <= 18'h14D06 ;
            12'd16 : y <= 18'h3E01B ;
            12'd17 : y <= 18'h14D06 ;
            12'd18 : y <= 18'h3E014 ;
            12'd19 : y <= 18'h2200A ;
            12'd20 : y <= 18'h20030 ;
            12'd21 : y <= 18'h09E00 ;
            12'd22 : y <= 18'h0DE10 ;
            12'd23 : y <= 18'h3A00A ;
            12'd24 : y <= 18'h01E00 ;
            12'd25 : y <= 18'h2FE00 ;
            12'd26 : y <= 18'h2200A ;
            12'd27 : y <= 18'h20030 ;
            12'd28 : y <= 18'h09E00 ;
            12'd29 : y <= 18'h0DE20 ;
            12'd30 : y <= 18'h3A00A ;
            12'd31 : y <= 18'h01E01 ;
            12'd32 : y <= 18'h2FE00 ;
            12'd33 : y <= 18'h2200A ;
            12'd34 : y <= 18'h20030 ;
            12'd35 : y <= 18'h09E00 ;
            12'd36 : y <= 18'h0DE40 ;
            12'd37 : y <= 18'h3A00A ;
            12'd38 : y <= 18'h01E02 ;
            12'd39 : y <= 18'h2FE00 ;
            12'd40 : y <= 18'h2200A ;
            12'd41 : y <= 18'h20030 ;
            12'd42 : y <= 18'h09E00 ;
            12'd43 : y <= 18'h0DE80 ;
            12'd44 : y <= 18'h3A00A ;
            12'd45 : y <= 18'h01E03 ;
            12'd46 : y <= 18'h2FE00 ;
            12'd47 : y <= 18'h2200A ;
            12'd48 : y <= 18'h01200 ;
            12'd49 : y <= 18'h0112E ;
            12'd50 : y <= 18'h010E0 ;
            12'd51 : y <= 18'h22038 ;
            12'd52 : y <= 18'h01203 ;
            12'd53 : y <= 18'h011A9 ;
            12'd54 : y <= 18'h01080 ;
            12'd55 : y <= 18'h22038 ;
            12'd56 : y <= 18'h00000 ;
            12'd57 : y <= 18'h19001 ;
            12'd58 : y <= 18'h1B100 ;
            12'd59 : y <= 18'h1B200 ;
            12'd60 : y <= 18'h36038 ;
            12'd61 : y <= 18'h25000 ;
            12'd62 : y <= 18'h0BC00 ;
            12'd63 : y <= 18'h11C01 ;
            12'd64 : y <= 18'h00BC0 ;
            12'd65 : y <= 18'h03B0F ;
            12'd66 : y <= 18'h1DB0A ;
            12'd67 : y <= 18'h3604A ;
            12'd68 : y <= 18'h11C06 ;
            12'd69 : y <= 18'h00BC0 ;
            12'd70 : y <= 18'h03BF0 ;
            12'd71 : y <= 18'h1DBA0 ;
            12'd72 : y <= 18'h3604A ;
            12'd73 : y <= 18'h01C00 ;
            12'd74 : y <= 18'h2DC00 ;
            12'd75 : y <= 18'h2FC00 ;
            12'd76 : y <= 18'h25000 ;
            12'd77 : y <= 18'h0BA01 ;
            12'd78 : y <= 18'h14A0C ;
            12'd79 : y <= 18'h2DA01 ;
            12'd80 : y <= 18'h2FA01 ;
            12'd81 : y <= 18'h25000 ;
            12'd82 : y <= 18'h00000 ;
            12'd83 : y <= 18'h00000 ;
            12'd84 : y <= 18'h28000 ;
            12'd85 : y <= 18'h2004D ;
            12'd86 : y <= 18'h2003E ;
            12'd87 : y <= 18'h29001 ;
            12'd88 : y <= 18'h00000 ;
            12'd89 : y <= 18'h00000 ;
            default : y <= 18'd0 ;
       endcase
    end
end
endmodule 
